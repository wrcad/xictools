Josephson junctions I-V curve demo

*
* One can plot a pretty decent iv curve using transient analysis.
* This will show the differences between the various model options.
*
b1 1 0 phase jjva 
v1 2 0 pwl(0 0 2n 700m 4n 0 5n 0  7n -700m 9n 0)
r1 2 1 500
.model jjva b(level=2 mfactor=0.3)
 
.control
tran 5p 10n
plot -v1#branch vs v(1)
.endc

