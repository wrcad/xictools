* Josephson Interferometer demo
*
* This is a symmetric two junction interferometer.
*
* the squid loop
b1 1 0 100 jj1
b2 3 0 101 jj1
l1 1 2 2pH
l2 2 3 2pH
*
* the coupled control line
l3 4 5 2pH
l4 5 0 2pH
k1 l1 l3 .98
k2 l2 l4 .98
*
* damping resistance
rd1 1 0 .50
rd2 3 0 .50
*rd1 1 0 2
*rd2 3 0 2
*
* gate power supply
rg 2 10 50
vg 10 0 pulse(0 80m 0p 20p)
*
* source power supply
rc 4 11 50
vc 11 0 pulse(0 25m 0 200p)
*vc 11 0 pulse(0 25.4m 50p 2p 2p)
*
.tran 1p 200p
*
* Type "run", then "plot v(11) v(3)" to display the control
* voltage and gate voltage.
*
* Initially, we have a single vortex transition.
*
* Suggestions for experiment:
*    1. raise the values of rd1 and rd2 and note the effects,
*    1. change the amplitude of vg, find the critical point,
*    3. change vc to a pulse source:
*       vc 11 0 pulse(0 50m 50p 2p 2p)
*       and find the amplitude where switching is metastable
*
*Nb 2500 A/cm2   area = 40 square microns
.model jj1 jj(rtype=1,cct=1,icon=10m,vg=2.8m,delv=0.08m,
+ icrit=1m,r0=30,rn=1.647059,cap=1.548944p)
.end

.control
run
plot v(11) v(1) ysep
edit
.endc
