* Josephson flux shuttle shift register operating range analysis\n\n\
To run, give these commands to WRspice after sourcing this file:\n\
    mplot -on\n\
    check
*
*
* Warning:  This file probably requires WRspice-4.3.3 or later.
* Warning:  This uses WRspice extensions, file is not portable.
* 
.check

* Set this to 0 to use TRAN ramp-up and uic instead of DCOP.
.param dcop=1

* Below,
* Level=1 selects the internal RSJ JJ model.
* Level=2 selects the example Verilog-A JJ model, if loaded (with
* the devload command).
* Level=3 selects the internal microscopic JJ model.
*
.model jj1 jj(level=1)

.if dcop
.tran 1p 400p
.else
.tran 1p 400p uic
.endif

.exec
# Margins of a Josephson flux shuttle shift register
# This is an example of an operating range analysis input file
#
compose checkPNTS values 61p 101p 141p 181p 221p 261p 301p
checkFAIL = 0
# above two lines are required in header, the rest are optional
#
# central value of first variable, number of evaluation steps above and
# below, step delta:
checkVAL1 = .4
checkSTP1 = 3
checkDEL1 = .1
#
# same thing for second variable
checkVAL2 = 120
checkSTP2 = 3
checkDEL2 = 10
#
# end of header
.endc
.control
#
# The following code is evaluated just after the time variable exceeds
# each one of the checkPNTS
#
if time > checkPNTS[0]
        if time < checkPNTS[1]
                checkFAIL = 0
                if abs(v(100) - v(101) - 5.3) > 2
                        checkFAIL = 1;
                end
                if abs(v(101) - v(102)) > 2
                        checkFAIL = 1;
                end
                if abs(v(102) - v(103)) > 2
                        checkFAIL = 1;
                end
                if abs(v(103) - v(104)) > 2
                        checkFAIL = 1;
                end
                if abs(v(104) - v(105)) > 2
                        checkFAIL = 1;
                end
                if abs(v(105) - v(106)) > 2
                        checkFAIL = 1;
                end
                echo tp1
        end
end
if time > checkPNTS[1]
        if time < checkPNTS[2]
                checkFAIL = 0
                if abs(v(100) - v(101)) > 2
                        checkFAIL = 1;
                end
                if abs(v(101) - v(102) - 5.3) > 2
                        checkFAIL = 1;
                end
                if abs(v(102) - v(103)) > 2
                        checkFAIL = 1;
                end
                if abs(v(103) - v(104)) > 2
                        checkFAIL = 1;
                end
                if abs(v(104) - v(105)) > 2
                        checkFAIL = 1;
                end
                if abs(v(105) - v(106)) > 2
                        checkFAIL = 1;
                end
                echo tp2
        end
end
if time > checkPNTS[2]
        if time < checkPNTS[3]
                checkFAIL = 0
                if abs(v(100) - v(101)) > 2
                        checkFAIL = 1;
                end
                if abs(v(101) - v(102)) > 2
                        checkFAIL = 1;
                end
                if abs(v(102) - v(103) - 5.3) > 2
                        checkFAIL = 1;
                end
                if abs(v(103) - v(104)) > 2
                        checkFAIL = 1;
                end
                if abs(v(104) - v(105)) > 2
                        checkFAIL = 1;
                end
                if abs(v(105) - v(106)) > 2
                        checkFAIL = 1;
                end
                echo tp3
        end
end
if time > checkPNTS[3]
        if time < checkPNTS[4]
                checkFAIL = 0
                if abs(v(100) - v(101)) > 2
                        checkFAIL = 1;
                end
                if abs(v(101) - v(102)) > 2
                        checkFAIL = 1;
                end
                if abs(v(102) - v(103)) > 2
                        checkFAIL = 1;
                end
                if abs(v(103) - v(104) - 5.3) > 2
                        checkFAIL = 1;
                end
                if abs(v(104) - v(105)) > 2
                        checkFAIL = 1;
                end
                if abs(v(105) - v(106)) > 2
                        checkFAIL = 1;
                end
                echo tp4
        end
end
if time > checkPNTS[4]
        if time < checkPNTS[5]
                checkFAIL = 0
                if abs(v(100) - v(101)) > 2
                        checkFAIL = 1;
                end
                if abs(v(101) - v(102)) > 2
                        checkFAIL = 1;
                end
                if abs(v(102) - v(103)) > 2
                        checkFAIL = 1;
                end
                if abs(v(103) - v(104)) > 2
                        checkFAIL = 1;
                end
                if abs(v(104) - v(105) - 5.3) > 2
                        checkFAIL = 1;
                end
                if abs(v(105) - v(106)) > 2
                        checkFAIL = 1;
                end
                echo tp5
        end
end
if time > checkPNTS[5]
        if time < checkPNTS[6]
                checkFAIL = 0
                if abs(v(100) - v(101)) > 2
                        checkFAIL = 1;
                end
                if abs(v(101) - v(102)) > 2
                        checkFAIL = 1;
                end
                if abs(v(102) - v(103)) > 2
                        checkFAIL = 1;
                end
                if abs(v(103) - v(104)) > 2
                        checkFAIL = 1;
                end
                if abs(v(104) - v(105)) > 2
                        checkFAIL = 1;
                end
                if abs(v(105) - v(106) - 5.3) > 2
                        checkFAIL = 1;
                end
                echo tp6
        end
end
if time > checkPNTS[6]
        checkFAIL = 0
        if abs(v(100) - v(101)) > 2
                checkFAIL = 1;
        end
        if abs(v(101) - v(102)) > 2
                checkFAIL = 1;
        end
        if abs(v(102) - v(103)) > 2
                checkFAIL = 1;
        end
        if abs(v(103) - v(104)) > 2
                checkFAIL = 1;
        end
        if abs(v(104) - v(105)) > 2
                checkFAIL = 1;
        end
        if abs(v(105) - v(106)) > 2
                checkFAIL = 1;
        end
end
.endc

r1 1 2 100
r2 2 0 $value1
r3 3 0 $value1
r4 4 0 $value1
r5 5 0 $value1
r6 6 0 $value1
r7 7 0 $value1
r8 8 0 $value1
r9 9 0 $value1
r10 10 11 100
r20 20 21 100
r30 30 31 100

l1 2 3 3p
l2 3 4 3p
l3 4 5 3p
l4 5 6 3p
l5 6 7 3p
l6 7 8 3p
l7 8 9 3p

l10 11 12 3p
l11 12 13 3p
l12 13 0  3p
l20 21 22 3p
l21 22 0  3p
l30 31 32 3p
l31 32 0  3p

k1 l10 l1 .99
k2 l11 l4 .99
k3 l12 l7 .99
k4 l20 l2 .99
k5 l21 l5 .99
k6 l30 l3 .99
k7 l31 l6 .99

b1 2 0 100 jj1
b2 3 0 101 jj1
b3 4 0 102 jj1
b4 5 0 103 jj1
b5 6 0 104 jj1
b6 7 0 105 jj1
b7 8 0 106 jj1
b8 9 0 107 jj1

* Three-phase clock
v1 10 0 pulse(0 $value2%m   25p 10p 10p 10p 120p)
v2 20 0 pulse(0 $value2%m  65p 10p 10p 10p 120p)
v3 30 0 pulse(0 $value2%m 105p 10p 10p 10p 120p)

v4 1 0 pulse(0 40m 25p 10p 10p)

