module integer_example;

integer counter; // general purpose variable used as a counter.
initial
	counter = -1; // A negative one is stored in the counter

endmodule


