* \nExample parameter range analysis of NOR gate.

* We need to save the special vectors accessed for pass/fail testing.
.save @b2.x3[n]
.save @b3.x3[n]

.tran 0.1p 1n

* This is called periodically during simulation, performs pass/fail test.
.control cb

  # Compare expected result to analog, quit if different.
  if ($&v(102) eq $&(@B2.X3[n]-@B3.X3[n]))
#    echo ERROR time=$&time : $&v(102) $&(@B2.X3[n]-@B3.X3[n])
    return 0
  end
  return 1
.endc

* Logical result for comparison in pass/fail test.
vout 102 0 pulse(0 1 DLY+2*PER-10p 0.2p 0.2p 0.5*PER-0.2p PER BD1) |
+ pulse(0 1 DLY+2*PER-10p 0.2p 0.2p 0.5*PER-0.2p PER BD2)

.control

# First do a run and plot the results.  This is not needed and the
# following two lines can be commented.
#run
#plot ysep v(3) v(6) v(8) v(5) v(15) v(102) (@b2.x3[n]-@b3.x3[n])

# Enable operating point limit search to depth.
set checkiterate=6

# Unbind any "control" codeblock (unlikely to be one).  Since we call
# check from the .control block here, the .control block will not be
# bound as it would be in a normal operating range input file.
codeblock -b

# Start incremental margin analysis.
check -b

# Below, find the operating range of the circuit parameters listed. 
# The second findrange argument is quoted so it is taken as a name
# string and not parameter expanded, as it is in the final argument.

# Some of these may generate warning messages as the search takes
# parameters out of range.  Some parameters may not have an upper or
# lower bound.

findrange -n1 "b0ics" b0.x0,ics b0ics
echo b0.x0 ics
print b0ics_min b0ics_max 0.5*(b0ics_min+b0ics_max)  b0ics

findrange -n1 "b1ics" b1.x0,ics b1ics
echo b1.x0 ics
print b1ics_min b1ics_max 0.5*(b1ics_min+b1ics_max)  b1ics

findrange -n1 "b2ics" b2.x0,ics b2ics
echo b2.x0 ics
print b2ics_min b2ics_max 0.5*(b2ics_min+b2ics_max)  b2ics

findrange -n1 "b3ics" b3.x0,ics b3ics
echo b3.x0 ics
print b3ics_min b3ics_max 0.5*(b3ics_min+b3ics_max)  b3ics

findrange -n1 "b4ics" b4.x0,ics b4ics
echo b4.x0 ics
print b4ics_min b4ics_max 0.5*(b4ics_min+b4ics_max)  b4ics

findrange -n1 "b5ics" b5.x0,ics b5ics
echo b5.x0 ics
print b5ics_min b5ics_max 0.5*(b5ics_min+b5ics_max)  b5ics

findrange -n1 "b6ics" b6.x0,ics b6ics
echo b6.x0 ics
print b6ics_min b6ics_max 0.5*(b6ics_min+b6ics_max)  b6ics

findrange -n1 "b7ics" b7.x0,ics b7ics
echo b7.x0 ics
print b7ics_min b7ics_max 0.5*(b7ics_min+b7ics_max)  b7ics

findrange -n1 "r0r" r0.x0,r r0r
echo r0.x0 r
print r0r_min r0r_max 0.5*(r0r_min+r0r_max)  r0r

findrange -n1 "r1r" r1.x0,r r1r
echo r1.x0 r
print r1r_min r1r_max 0.5*(r1r_min+r1r_max)  r1r

findrange -n1 "r2r" r2.x0,r r2r
echo r2.x0 r
print r2r_min r2r_max 0.5*(r2r_min+r2r_max)  r2r

findrange -n1 "r3r" r3.x0,r r3r
echo r3.x0 r
print r3r_min r3r_max 0.5*(r3r_min+r3r_max)  r0r

findrange -n1 "l5l" l5.x0,l l5l
echo l5.x0 l
print l5l_min l5l_max 0.5*(l5l_min+l5l_max)  l5l

# End the incremental range analysis.
check -c

.endc

* Set up periodic result checking (call cb periodically).
.stop tran at DLY+PER repeat PER call cb silent

* Set up run parameters, input patterns are included here in this example.
.param BD1="bprbs6 r=-1"
.param BD2="bprbs6 rb=11 r=-1"
.param PER=50pS
.param DLY=20pS

* Nominal values of parameters to be varied.
.param b0ics=140u
.param b1ics=250u
.param b2ics=310u
.param b3ics=174u
.param b4ics=294u
.param b5ics=355u
.param b6ics=294u
.param b7ics=264u
.param r0r=40
.param r1r=42
.param r2r=74
.param r3r=65
.param l5l=5.88p

* The circuit:  a NOR gate created from the rsfq_lib library.
* Generated by Xic from cell nor_test
*.tran 0.1p 1n
*.plot tran v(3) v(6) v(8) v(5) v(15)
.model jj5ee jj(VSHUNT=0.6857mV)
LT0 2 12 3.3p
LT1 9 13 3.3p
LT2 10 14 3.3p
V0 2 0 gpulse(0 0 DLY+15p 2p PER BD1)
V1 9 0 gpulse(0 0 DLY+10p 2p PER BD2)
V2 10 0 gpulse(0 0 DLY 2p PER)
V3 VDD 0 10m
X0 4 8 5 VDD inv
X1 12 3 VDD jtl
X2 3 6 4 VDD conf_il
X3 5 15 7 VDD dff
X4 13 6 VDD jtl
X5 11 8 7 VDD split
X6 14 11 VDD jtl
.subckt inv 26 27 28 VBIAS
B0 10 11 29 jj5ee ics=b0ics
B1 9 15 30  jj5ee ics=b1ics
B2 10 16 31 jj5ee ics=b2ics
B3 12 17 32 jj5ee ics=b3ics
B4 13 18 33 jj5ee ics=b4ics
B5 14 19 34 jj5ee ics=b5ics
B6 21 24 35 jj5ee ics=b6ics
B7 23 25 36 jj5ee ics=b7ics
L0 26 9 2pH
L1 9 6 1.03pH
L2 6 10 .97pH
L3 11 12 .97pH
L4 12 7 .33pH
L5 7 13 l5l
L6 8 13 1.3pH
L7 14 8 1.02pH
L8 27 14 .79pH
L9 17 20 1.04pH
L10 20 18 .57pH
L11 20 21 .875pH
L12 21 22 1.7pH
L13 22 23 1.11pH
L14 23 28 2.37pH
LP0 3 6 .35pH
LP1 4 7 .57pH
LP2 5 8 .33pH
LP3 15 0 .03pH
LP4 16 0 .09pH
LP5 19 0 .02pH
LP6 2 22 .5pH
LP7 24 0 .145pH
LP8 25 0 .03pH
R0 VBIAS 3 r0r
R1 VBIAS 4 r1r
R2 VBIAS 5 r2r
R3 VBIAS 2 r3r
.ends inv
.subckt jtl IN OUT VBIAS
B0 5 7 9 jj5ee ics=250u
B1 6 8 10 jj5ee ics=250u
LP0 7 0 .1pH
LP1 8 0 .1pH
LT0 IN 5 2.1pH
LT1 5 4 2.1pH
LT2 4 6 2.1pH
LT3 6 OUT 2.1pH
R0 VBIAS 4 29
.ends jtl
.subckt conf_il IN1 IN2 OUT VBIAS
B0 8 7 15 jj5ee ics=350u
B1 8 9 16 jj5ee ics=200u
B2 11 10 17 jj5ee ics=200u
B3 11 13 18 jj5ee ics=350u
B4 12 14 19 jj5ee ics=300u
LP0 7 0 0.25pH
LP1 13 0 0.25pH
LP2 14 0 0.26pH
LT0 IN1 8 1.87pH
LT1 9 5 1.39pH
LT2 IN2 11 1.87pH
LT3 10 5 1.39pH
LT4 5 6 0.44pH
LT5 6 12 1.94pH
LT6 12 OUT 1.80pH
R0 VBIAS 6 18
.ends conf_il
.subckt dff IN OUT CLK VBIAS
B0 6 7 9 jj5ee ics=270u
B1 8 5 10 jj5ee ics=245u
B2 5 0 11 jj5ee ics=245u
B3 7 0 12 jj5ee ics=270u
L0 5 7 8.46pH
LT0 CLK 6 1.58pH
LT1 IN 8 2.76pH
LT2 7 OUT 3.16pH
R0 VBIAS 5 59
.ends dff
.subckt split IN OUT1 OUT2 VBIAS
B0 9 7 14 jj5ee ics=250u
B1 10 11 15 jj5ee ics=355u
B2 12 13 16 jj5ee ics=250u
LP0 7 0 0.05pH
LP1 8 6 0.13pH
LP2 11 0 0.05pH
LP3 13 0 0.05pH
LT0 5 9 1.63pH
LT1 9 OUT2 1.98pH
LT2 IN 10 0.82pH
LT3 10 6 1.16pH
LT4 6 5 0.05pH
LT5 5 12 1.63pH
LT6 12 OUT1 1.98pH
R0 VBIAS 8 17
.ends split

