
module time_example;

time save_sim_time; // Define a time variable save_sim_time
initial
	save_sim_time = $time; // Save the current simulation time 

endmodule
