/****************************************************************************
 *                                                                          *
 *  VERILOG HIGH-LEVEL DESCRIPTION OF THE ISCAS-85 BENCHMARK CIRCUIT c6288  *
 *                                                                          *
 *  Function: 16 x 16 Multiplier                                            *
 *                                                                          *
 *  Written by: Mark C. Hansen                                              *
 *                                                                          *
 *  Last modified: Nov 12, 1997                                             *
 *                                                                          *
 ****************************************************************************/

module m16x16 (in256, in239, in222, in205, in188, in171, in154, in137, 
                 in120, in103, in86, in69, in52, in35, in18, in1,
                 in528, in511, in494, in477, in460, in443, in426, in409,
                 in392, in375, in358, in341, in324, in307, in290, in273,
                 out6287, out6288, out6280, out6270,
                 out6260, out6250, out6240, out6230, 
                 out6220, out6210, out6200, out6190, 
                 out6180, out6170, out6160, out6150, 
                 out6123, out5971, out5672, out5308, 
                 out4946, out4591, out4241, out3895,
                 out3552, out3211, out2877, out2548,
                 out2223, out1901, out1581, out545);

  input          in256, in239, in222, in205, in188, in171, in154, in137, 
                 in120, in103, in86, in69, in52, in35, in18, in1,
                 in528, in511, in494, in477, in460, in443, in426, in409,
                 in392, in375, in358, in341, in324, in307, in290, in273;
  output         out6287, out6288, out6280, out6270,
                 out6260, out6250, out6240, out6230, 
                 out6220, out6210, out6200, out6190, 
                 out6180, out6170, out6160, out6150, 
                 out6123, out5971, out5672, out5308, 
                 out4946, out4591, out4241, out3895,
                 out3552, out3211, out2877, out2548,
                 out2223, out1901, out1581, out545;

  reg [15:0]   A, B;
  wire [31:0]   P,P1,P2;

  initial 
    begin
      # 1;
      A = 0101010101010101; B= 1111_1111_1111_1111;
      # 1;
      $display("A=%h,B=%h,P=%h,P1=%h,P2=%h",A,B,P,P1,P2);
      A = 1010101010101010; B= 1111111111111111;
      # 1;
      $display("A=%h,B=%h,P=%h,P1=%h,P2=%h",A,B,P,P1,P2);
      A = 0101010101010101; B= 1101111111111111;
      # 1;
      $display("A=%h,B=%h,P=%h,P1=%h,P2=%h",A,B,P,P1,P2);
      A = 1010101010101010; B= 1101111111111111;
      # 1;
      $display("A=%h,B=%h,P=%h,P1=%h,P2=%h",A,B,P,P1,P2);
      A = 1101101101101101; B= 1111111111111111;
      # 1;
      $display("A=%h,B=%h,P=%h,P1=%h,P2=%h",A,B,P,P1,P2);
      A = 0110110110110110; B= 1111111111111111;
      # 1;
      $display("A=%h,B=%h,P=%h,P1=%h,P2=%h",A,B,P,P1,P2);
      A = 1011011011011011; B= 1111111111111111;
      # 1;
      $display("A=%h,B=%h,P=%h,P1=%h,P2=%h",A,B,P,P1,P2);
      A = 1111111111111111; B= 1101010101010101;
      # 1;
      $display("A=%h,B=%h,P=%h,P1=%h,P2=%h",A,B,P,P1,P2);
      A = 1111111111111111; B= 0110101010101010;
      # 1;
      $display("A=%h,B=%h,P=%h,P1=%h,P2=%h",A,B,P,P1,P2);
      A = 1111111111111110; B= 1101010101010101;
      # 1;
      $display("A=%h,B=%h,P=%h,P1=%h,P2=%h",A,B,P,P1,P2);
      A = 1111111111111110; B= 0110101010101010;
      # 1;
      $display("A=%h,B=%h,P=%h,P1=%h,P2=%h",A,B,P,P1,P2);
      A = 1111111111111111; B= 0000000000000000;
      # 1;
      $display("A=%h,B=%h,P=%h,P1=%h,P2=%h",A,B,P,P1,P2);
    end
	
  TopLevel6288 Ckt6288 (A, B, P);
  TopLevel6288 Ckt6288_a (A, P[15:0], P1);
  TopLevel6288 Ckt6288_b (B, P[15:0], P2);

endmodule /* Circuit6288 */

/*************************************************************************/

module TopLevel6288 (A, B, P);

  input[15:0]	A, B;
  output[31:0]	P;

  wire          C14_15, S14_15, S13_15, S12_15,
               S11_15, S10_15, S9_15, S8_15,
               S7_15, S6_15, S5_15, S4_15,
               S3_15, S2_15, S1_15, S0_15,
               S0_14, S0_13, S0_12, S0_11,
               S0_10, S0_9, S0_8, S0_7,
               S0_6, S0_5, S0_4, S0_3,
               S0_2, S0_1, S0_0, A0B0;

  assign
    P[31:0] = {C14_15, S14_15, S13_15, S12_15,
               S11_15, S10_15, S9_15, S8_15,
               S7_15, S6_15, S5_15, S4_15,
               S3_15, S2_15, S1_15, S0_15,
               S0_14, S0_13, S0_12, S0_11,
               S0_10, S0_9, S0_8, S0_7,
               S0_6, S0_5, S0_4, S0_3,
               S0_2, S0_1, S0_0, A0B0};

  and GA0B0(A0B0, A[0], B[0]);
  and GA0B1(A0B1, A[0], B[1]);
  and GA0B2(A0B2, A[0], B[2]);
  and GA0B3(A0B3, A[0], B[3]);
  and GA0B4(A0B4, A[0], B[4]);
  and GA0B5(A0B5, A[0], B[5]);
  and GA0B6(A0B6, A[0], B[6]);
  and GA0B7(A0B7, A[0], B[7]);
  and GA0B8(A0B8, A[0], B[8]);
  and GA0B9(A0B9, A[0], B[9]);
  and GA0B10(A0B10, A[0], B[10]);
  and GA0B11(A0B11, A[0], B[11]);
  and GA0B12(A0B12, A[0], B[12]);
  and GA0B13(A0B13, A[0], B[13]);
  and GA0B14(A0B14, A[0], B[14]);
  and GA0B15(A0B15, A[0], B[15]);

  and GA1B0(A1B0, A[1], B[0]);
  and GA1B1(A1B1, A[1], B[1]);
  and GA1B2(A1B2, A[1], B[2]);
  and GA1B3(A1B3, A[1], B[3]);
  and GA1B4(A1B4, A[1], B[4]);
  and GA1B5(A1B5, A[1], B[5]);
  and GA1B6(A1B6, A[1], B[6]);
  and GA1B7(A1B7, A[1], B[7]);
  and GA1B8(A1B8, A[1], B[8]);
  and GA1B9(A1B9, A[1], B[9]);
  and GA1B10(A1B10, A[1], B[10]);
  and GA1B11(A1B11, A[1], B[11]);
  and GA1B12(A1B12, A[1], B[12]);
  and GA1B13(A1B13, A[1], B[13]);
  and GA1B14(A1B14, A[1], B[14]);
  and GA1B15(A1B15, A[1], B[15]);

  and GA2B0(A2B0, A[2], B[0]);
  and GA2B1(A2B1, A[2], B[1]);
  and GA2B2(A2B2, A[2], B[2]);
  and GA2B3(A2B3, A[2], B[3]);
  and GA2B4(A2B4, A[2], B[4]);
  and GA2B5(A2B5, A[2], B[5]);
  and GA2B6(A2B6, A[2], B[6]);
  and GA2B7(A2B7, A[2], B[7]);
  and GA2B8(A2B8, A[2], B[8]);
  and GA2B9(A2B9, A[2], B[9]);
  and GA2B10(A2B10, A[2], B[10]);
  and GA2B11(A2B11, A[2], B[11]);
  and GA2B12(A2B12, A[2], B[12]);
  and GA2B13(A2B13, A[2], B[13]);
  and GA2B14(A2B14, A[2], B[14]);
  and GA2B15(A2B15, A[2], B[15]);

  and GA3B0(A3B0, A[3], B[0]);
  and GA3B1(A3B1, A[3], B[1]);
  and GA3B2(A3B2, A[3], B[2]);
  and GA3B3(A3B3, A[3], B[3]);
  and GA3B4(A3B4, A[3], B[4]);
  and GA3B5(A3B5, A[3], B[5]);
  and GA3B6(A3B6, A[3], B[6]);
  and GA3B7(A3B7, A[3], B[7]);
  and GA3B8(A3B8, A[3], B[8]);
  and GA3B9(A3B9, A[3], B[9]);
  and GA3B10(A3B10, A[3], B[10]);
  and GA3B11(A3B11, A[3], B[11]);
  and GA3B12(A3B12, A[3], B[12]);
  and GA3B13(A3B13, A[3], B[13]);
  and GA3B14(A3B14, A[3], B[14]);
  and GA3B15(A3B15, A[3], B[15]);

  and GA4B0(A4B0, A[4], B[0]);
  and GA4B1(A4B1, A[4], B[1]);
  and GA4B2(A4B2, A[4], B[2]);
  and GA4B3(A4B3, A[4], B[3]);
  and GA4B4(A4B4, A[4], B[4]);
  and GA4B5(A4B5, A[4], B[5]);
  and GA4B6(A4B6, A[4], B[6]);
  and GA4B7(A4B7, A[4], B[7]);
  and GA4B8(A4B8, A[4], B[8]);
  and GA4B9(A4B9, A[4], B[9]);
  and GA4B10(A4B10, A[4], B[10]);
  and GA4B11(A4B11, A[4], B[11]);
  and GA4B12(A4B12, A[4], B[12]);
  and GA4B13(A4B13, A[4], B[13]);
  and GA4B14(A4B14, A[4], B[14]);
  and GA4B15(A4B15, A[4], B[15]);

  and GA5B0(A5B0, A[5], B[0]);
  and GA5B1(A5B1, A[5], B[1]);
  and GA5B2(A5B2, A[5], B[2]);
  and GA5B3(A5B3, A[5], B[3]);
  and GA5B4(A5B4, A[5], B[4]);
  and GA5B5(A5B5, A[5], B[5]);
  and GA5B6(A5B6, A[5], B[6]);
  and GA5B7(A5B7, A[5], B[7]);
  and GA5B8(A5B8, A[5], B[8]);
  and GA5B9(A5B9, A[5], B[9]);
  and GA5B10(A5B10, A[5], B[10]);
  and GA5B11(A5B11, A[5], B[11]);
  and GA5B12(A5B12, A[5], B[12]);
  and GA5B13(A5B13, A[5], B[13]);
  and GA5B14(A5B14, A[5], B[14]);
  and GA5B15(A5B15, A[5], B[15]);

  and GA6B0(A6B0, A[6], B[0]);
  and GA6B1(A6B1, A[6], B[1]);
  and GA6B2(A6B2, A[6], B[2]);
  and GA6B3(A6B3, A[6], B[3]);
  and GA6B4(A6B4, A[6], B[4]);
  and GA6B5(A6B5, A[6], B[5]);
  and GA6B6(A6B6, A[6], B[6]);
  and GA6B7(A6B7, A[6], B[7]);
  and GA6B8(A6B8, A[6], B[8]);
  and GA6B9(A6B9, A[6], B[9]);
  and GA6B10(A6B10, A[6], B[10]);
  and GA6B11(A6B11, A[6], B[11]);
  and GA6B12(A6B12, A[6], B[12]);
  and GA6B13(A6B13, A[6], B[13]);
  and GA6B14(A6B14, A[6], B[14]);
  and GA6B15(A6B15, A[6], B[15]);

  and GA7B0(A7B0, A[7], B[0]);
  and GA7B1(A7B1, A[7], B[1]);
  and GA7B2(A7B2, A[7], B[2]);
  and GA7B3(A7B3, A[7], B[3]);
  and GA7B4(A7B4, A[7], B[4]);
  and GA7B5(A7B5, A[7], B[5]);
  and GA7B6(A7B6, A[7], B[6]);
  and GA7B7(A7B7, A[7], B[7]);
  and GA7B8(A7B8, A[7], B[8]);
  and GA7B9(A7B9, A[7], B[9]);
  and GA7B10(A7B10, A[7], B[10]);
  and GA7B11(A7B11, A[7], B[11]);
  and GA7B12(A7B12, A[7], B[12]);
  and GA7B13(A7B13, A[7], B[13]);
  and GA7B14(A7B14, A[7], B[14]);
  and GA7B15(A7B15, A[7], B[15]);

  and GA8B0(A8B0, A[8], B[0]);
  and GA8B1(A8B1, A[8], B[1]);
  and GA8B2(A8B2, A[8], B[2]);
  and GA8B3(A8B3, A[8], B[3]);
  and GA8B4(A8B4, A[8], B[4]);
  and GA8B5(A8B5, A[8], B[5]);
  and GA8B6(A8B6, A[8], B[6]);
  and GA8B7(A8B7, A[8], B[7]);
  and GA8B8(A8B8, A[8], B[8]);
  and GA8B9(A8B9, A[8], B[9]);
  and GA8B10(A8B10, A[8], B[10]);
  and GA8B11(A8B11, A[8], B[11]);
  and GA8B12(A8B12, A[8], B[12]);
  and GA8B13(A8B13, A[8], B[13]);
  and GA8B14(A8B14, A[8], B[14]);
  and GA8B15(A8B15, A[8], B[15]);

  and GA9B0(A9B0, A[9], B[0]);
  and GA9B1(A9B1, A[9], B[1]);
  and GA9B2(A9B2, A[9], B[2]);
  and GA9B3(A9B3, A[9], B[3]);
  and GA9B4(A9B4, A[9], B[4]);
  and GA9B5(A9B5, A[9], B[5]);
  and GA9B6(A9B6, A[9], B[6]);
  and GA9B7(A9B7, A[9], B[7]);
  and GA9B8(A9B8, A[9], B[8]);
  and GA9B9(A9B9, A[9], B[9]);
  and GA9B10(A9B10, A[9], B[10]);
  and GA9B11(A9B11, A[9], B[11]);
  and GA9B12(A9B12, A[9], B[12]);
  and GA9B13(A9B13, A[9], B[13]);
  and GA9B14(A9B14, A[9], B[14]);
  and GA9B15(A9B15, A[9], B[15]);

  and GA10B0(A10B0, A[10], B[0]);
  and GA10B1(A10B1, A[10], B[1]);
  and GA10B2(A10B2, A[10], B[2]);
  and GA10B3(A10B3, A[10], B[3]);
  and GA10B4(A10B4, A[10], B[4]);
  and GA10B5(A10B5, A[10], B[5]);
  and GA10B6(A10B6, A[10], B[6]);
  and GA10B7(A10B7, A[10], B[7]);
  and GA10B8(A10B8, A[10], B[8]);
  and GA10B9(A10B9, A[10], B[9]);
  and GA10B10(A10B10, A[10], B[10]);
  and GA10B11(A10B11, A[10], B[11]);
  and GA10B12(A10B12, A[10], B[12]);
  and GA10B13(A10B13, A[10], B[13]);
  and GA10B14(A10B14, A[10], B[14]);
  and GA10B15(A10B15, A[10], B[15]);

  and GA11B0(A11B0, A[11], B[0]);
  and GA11B1(A11B1, A[11], B[1]);
  and GA11B2(A11B2, A[11], B[2]);
  and GA11B3(A11B3, A[11], B[3]);
  and GA11B4(A11B4, A[11], B[4]);
  and GA11B5(A11B5, A[11], B[5]);
  and GA11B6(A11B6, A[11], B[6]);
  and GA11B7(A11B7, A[11], B[7]);
  and GA11B8(A11B8, A[11], B[8]);
  and GA11B9(A11B9, A[11], B[9]);
  and GA11B10(A11B10, A[11], B[10]);
  and GA11B11(A11B11, A[11], B[11]);
  and GA11B12(A11B12, A[11], B[12]);
  and GA11B13(A11B13, A[11], B[13]);
  and GA11B14(A11B14, A[11], B[14]);
  and GA11B15(A11B15, A[11], B[15]);

  and GA12B0(A12B0, A[12], B[0]);
  and GA12B1(A12B1, A[12], B[1]);
  and GA12B2(A12B2, A[12], B[2]);
  and GA12B3(A12B3, A[12], B[3]);
  and GA12B4(A12B4, A[12], B[4]);
  and GA12B5(A12B5, A[12], B[5]);
  and GA12B6(A12B6, A[12], B[6]);
  and GA12B7(A12B7, A[12], B[7]);
  and GA12B8(A12B8, A[12], B[8]);
  and GA12B9(A12B9, A[12], B[9]);
  and GA12B10(A12B10, A[12], B[10]);
  and GA12B11(A12B11, A[12], B[11]);
  and GA12B12(A12B12, A[12], B[12]);
  and GA12B13(A12B13, A[12], B[13]);
  and GA12B14(A12B14, A[12], B[14]);
  and GA12B15(A12B15, A[12], B[15]);

  and GA13B0(A13B0, A[13], B[0]);
  and GA13B1(A13B1, A[13], B[1]);
  and GA13B2(A13B2, A[13], B[2]);
  and GA13B3(A13B3, A[13], B[3]);
  and GA13B4(A13B4, A[13], B[4]);
  and GA13B5(A13B5, A[13], B[5]);
  and GA13B6(A13B6, A[13], B[6]);
  and GA13B7(A13B7, A[13], B[7]);
  and GA13B8(A13B8, A[13], B[8]);
  and GA13B9(A13B9, A[13], B[9]);
  and GA13B10(A13B10, A[13], B[10]);
  and GA13B11(A13B11, A[13], B[11]);
  and GA13B12(A13B12, A[13], B[12]);
  and GA13B13(A13B13, A[13], B[13]);
  and GA13B14(A13B14, A[13], B[14]);
  and GA13B15(A13B15, A[13], B[15]);

  and GA14B0(A14B0, A[14], B[0]);
  and GA14B1(A14B1, A[14], B[1]);
  and GA14B2(A14B2, A[14], B[2]);
  and GA14B3(A14B3, A[14], B[3]);
  and GA14B4(A14B4, A[14], B[4]);
  and GA14B5(A14B5, A[14], B[5]);
  and GA14B6(A14B6, A[14], B[6]);
  and GA14B7(A14B7, A[14], B[7]);
  and GA14B8(A14B8, A[14], B[8]);
  and GA14B9(A14B9, A[14], B[9]);
  and GA14B10(A14B10, A[14], B[10]);
  and GA14B11(A14B11, A[14], B[11]);
  and GA14B12(A14B12, A[14], B[12]);
  and GA14B13(A14B13, A[14], B[13]);
  and GA14B14(A14B14, A[14], B[14]);
  and GA14B15(A14B15, A[14], B[15]);

  and GA15B0(A15B0, A[15], B[0]);
  and GA15B1(A15B1, A[15], B[1]);
  and GA15B2(A15B2, A[15], B[2]);
  and GA15B3(A15B3, A[15], B[3]);
  and GA15B4(A15B4, A[15], B[4]);
  and GA15B5(A15B5, A[15], B[5]);
  and GA15B6(A15B6, A[15], B[6]);
  and GA15B7(A15B7, A[15], B[7]);
  and GA15B8(A15B8, A[15], B[8]);
  and GA15B9(A15B9, A[15], B[9]);
  and GA15B10(A15B10, A[15], B[10]);
  and GA15B11(A15B11, A[15], B[11]);
  and GA15B12(A15B12, A[15], B[12]);
  and GA15B13(A15B13, A[15], B[13]);
  and GA15B14(A15B14, A[15], B[14]);
  and GA15B15(A15B15, A[15], B[15]);

/* HA MHA0_0(S0_0,C0_0,A1B0,A0B1); */
not gn1_0_0(n1_0_0, A1B0);
not gn2_0_0(n2_0_0, n1_0_0);
nor gn3_0_0(n3_0_0, A1B0, n1_0_0);
nor gn4_0_0(n4_0_0, n2_0_0, n3_0_0);
nor gn5_0_0(n5_0_0, A0B1, n4_0_0);
nor gn6_0_0(n6_0_0, A0B1, n5_0_0);
nor gn7_0_0(n7_0_0, n4_0_0, n5_0_0);
nor gn8_0_0(S0_0, n6_0_0, n7_0_0);
nor gn9_0_0(C0_0, n1_0_0, n5_0_0);

/* HA MHA1_0(S1_0,C1_0,A2B0,A1B1); */
not gn1_1_0(n1_1_0, A2B0);
not gn2_1_0(n2_1_0, n1_1_0);
nor gn3_1_0(n3_1_0, A2B0, n1_1_0);
nor gn4_1_0(n4_1_0, n2_1_0, n3_1_0);
nor gn5_1_0(n5_1_0, A1B1, n4_1_0);
nor gn6_1_0(n6_1_0, A1B1, n5_1_0);
nor gn7_1_0(n7_1_0, n4_1_0, n5_1_0);
nor gn8_1_0(S1_0, n6_1_0, n7_1_0);
nor gn9_1_0(C1_0, n1_1_0, n5_1_0);

/* HA MHA2_0(S2_0,C2_0,A3B0,A2B1); */
not gn1_2_0(n1_2_0, A3B0);
not gn2_2_0(n2_2_0, n1_2_0);
nor gn3_2_0(n3_2_0, A3B0, n1_2_0);
nor gn4_2_0(n4_2_0, n2_2_0, n3_2_0);
nor gn5_2_0(n5_2_0, A2B1, n4_2_0);
nor gn6_2_0(n6_2_0, A2B1, n5_2_0);
nor gn7_2_0(n7_2_0, n4_2_0, n5_2_0);
nor gn8_2_0(S2_0, n6_2_0, n7_2_0);
nor gn9_2_0(C2_0, n1_2_0, n5_2_0);

/* HA MHA3_0(S3_0,C3_0,A4B0,A3B1); */
not gn1_3_0(n1_3_0, A4B0);
not gn2_3_0(n2_3_0, n1_3_0);
nor gn3_3_0(n3_3_0, A4B0, n1_3_0);
nor gn4_3_0(n4_3_0, n2_3_0, n3_3_0);
nor gn5_3_0(n5_3_0, A3B1, n4_3_0);
nor gn6_3_0(n6_3_0, A3B1, n5_3_0);
nor gn7_3_0(n7_3_0, n4_3_0, n5_3_0);
nor gn8_3_0(S3_0, n6_3_0, n7_3_0);
nor gn9_3_0(C3_0, n1_3_0, n5_3_0);

/* HA MHA4_0(S4_0,C4_0,A5B0,A4B1); */
not gn1_4_0(n1_4_0, A5B0);
not gn2_4_0(n2_4_0, n1_4_0);
nor gn3_4_0(n3_4_0, A5B0, n1_4_0);
nor gn4_4_0(n4_4_0, n2_4_0, n3_4_0);
nor gn5_4_0(n5_4_0, A4B1, n4_4_0);
nor gn6_4_0(n6_4_0, A4B1, n5_4_0);
nor gn7_4_0(n7_4_0, n4_4_0, n5_4_0);
nor gn8_4_0(S4_0, n6_4_0, n7_4_0);
nor gn9_4_0(C4_0, n1_4_0, n5_4_0);

/* HA MHA5_0(S5_0,C5_0,A6B0,A5B1); */
not gn1_5_0(n1_5_0, A6B0);
not gn2_5_0(n2_5_0, n1_5_0);
nor gn3_5_0(n3_5_0, A6B0, n1_5_0);
nor gn4_5_0(n4_5_0, n2_5_0, n3_5_0);
nor gn5_5_0(n5_5_0, A5B1, n4_5_0);
nor gn6_5_0(n6_5_0, A5B1, n5_5_0);
nor gn7_5_0(n7_5_0, n4_5_0, n5_5_0);
nor gn8_5_0(S5_0, n6_5_0, n7_5_0);
nor gn9_5_0(C5_0, n1_5_0, n5_5_0);

/* HA MHA6_0(S6_0,C6_0,A7B0,A6B1); */
not gn1_6_0(n1_6_0, A7B0);
not gn2_6_0(n2_6_0, n1_6_0);
nor gn3_6_0(n3_6_0, A7B0, n1_6_0);
nor gn4_6_0(n4_6_0, n2_6_0, n3_6_0);
nor gn5_6_0(n5_6_0, A6B1, n4_6_0);
nor gn6_6_0(n6_6_0, A6B1, n5_6_0);
nor gn7_6_0(n7_6_0, n4_6_0, n5_6_0);
nor gn8_6_0(S6_0, n6_6_0, n7_6_0);
nor gn9_6_0(C6_0, n1_6_0, n5_6_0);

/* HA MHA7_0(S7_0,C7_0,A8B0,A7B1); */
not gn1_7_0(n1_7_0, A8B0);
not gn2_7_0(n2_7_0, n1_7_0);
nor gn3_7_0(n3_7_0, A8B0, n1_7_0);
nor gn4_7_0(n4_7_0, n2_7_0, n3_7_0);
nor gn5_7_0(n5_7_0, A7B1, n4_7_0);
nor gn6_7_0(n6_7_0, A7B1, n5_7_0);
nor gn7_7_0(n7_7_0, n4_7_0, n5_7_0);
nor gn8_7_0(S7_0, n6_7_0, n7_7_0);
nor gn9_7_0(C7_0, n1_7_0, n5_7_0);

/* HA MHA8_0(S8_0,C8_0,A9B0,A8B1); */
not gn1_8_0(n1_8_0, A9B0);
not gn2_8_0(n2_8_0, n1_8_0);
nor gn3_8_0(n3_8_0, A9B0, n1_8_0);
nor gn4_8_0(n4_8_0, n2_8_0, n3_8_0);
nor gn5_8_0(n5_8_0, A8B1, n4_8_0);
nor gn6_8_0(n6_8_0, A8B1, n5_8_0);
nor gn7_8_0(n7_8_0, n4_8_0, n5_8_0);
nor gn8_8_0(S8_0, n6_8_0, n7_8_0);
nor gn9_8_0(C8_0, n1_8_0, n5_8_0);

/* HA MHA9_0(S9_0,C9_0,A10B0,A9B1); */
not gn1_9_0(n1_9_0, A10B0);
not gn2_9_0(n2_9_0, n1_9_0);
nor gn3_9_0(n3_9_0, A10B0, n1_9_0);
nor gn4_9_0(n4_9_0, n2_9_0, n3_9_0);
nor gn5_9_0(n5_9_0, A9B1, n4_9_0);
nor gn6_9_0(n6_9_0, A9B1, n5_9_0);
nor gn7_9_0(n7_9_0, n4_9_0, n5_9_0);
nor gn8_9_0(S9_0, n6_9_0, n7_9_0);
nor gn9_9_0(C9_0, n1_9_0, n5_9_0);

/* HA MHA10_0(S10_0,C10_0,A11B0,A10B1); */
not gn1_10_0(n1_10_0, A11B0);
not gn2_10_0(n2_10_0, n1_10_0);
nor gn3_10_0(n3_10_0, A11B0, n1_10_0);
nor gn4_10_0(n4_10_0, n2_10_0, n3_10_0);
nor gn5_10_0(n5_10_0, A10B1, n4_10_0);
nor gn6_10_0(n6_10_0, A10B1, n5_10_0);
nor gn7_10_0(n7_10_0, n4_10_0, n5_10_0);
nor gn8_10_0(S10_0, n6_10_0, n7_10_0);
nor gn9_10_0(C10_0, n1_10_0, n5_10_0);

/* HA MHA11_0(S11_0,C11_0,A12B0,A11B1); */
not gn1_11_0(n1_11_0, A12B0);
not gn2_11_0(n2_11_0, n1_11_0);
nor gn3_11_0(n3_11_0, A12B0, n1_11_0);
nor gn4_11_0(n4_11_0, n2_11_0, n3_11_0);
nor gn5_11_0(n5_11_0, A11B1, n4_11_0);
nor gn6_11_0(n6_11_0, A11B1, n5_11_0);
nor gn7_11_0(n7_11_0, n4_11_0, n5_11_0);
nor gn8_11_0(S11_0, n6_11_0, n7_11_0);
nor gn9_11_0(C11_0, n1_11_0, n5_11_0);

/* HA MHA12_0(S12_0,C12_0,A13B0,A12B1); */
not gn1_12_0(n1_12_0, A13B0);
not gn2_12_0(n2_12_0, n1_12_0);
nor gn3_12_0(n3_12_0, A13B0, n1_12_0);
nor gn4_12_0(n4_12_0, n2_12_0, n3_12_0);
nor gn5_12_0(n5_12_0, A12B1, n4_12_0);
nor gn6_12_0(n6_12_0, A12B1, n5_12_0);
nor gn7_12_0(n7_12_0, n4_12_0, n5_12_0);
nor gn8_12_0(S12_0, n6_12_0, n7_12_0);
nor gn9_12_0(C12_0, n1_12_0, n5_12_0);

/* HA MHA13_0(S13_0,C13_0,A14B0,A13B1); */
not gn1_13_0(n1_13_0, A14B0);
not gn2_13_0(n2_13_0, n1_13_0);
nor gn3_13_0(n3_13_0, A14B0, n1_13_0);
nor gn4_13_0(n4_13_0, n2_13_0, n3_13_0);
nor gn5_13_0(n5_13_0, A13B1, n4_13_0);
nor gn6_13_0(n6_13_0, A13B1, n5_13_0);
nor gn7_13_0(n7_13_0, n4_13_0, n5_13_0);
nor gn8_13_0(S13_0, n6_13_0, n7_13_0);
nor gn9_13_0(C13_0, n1_13_0, n5_13_0);

/* HA MHA14_0(S14_0,C14_0,A15B0,A14B1); */
not gn1_14_0(n1_14_0, A15B0);
not gn2_14_0(n2_14_0, n1_14_0);
nor gn3_14_0(n3_14_0, A15B0, n1_14_0);
nor gn4_14_0(n4_14_0, n2_14_0, n3_14_0);
nor gn5_14_0(n5_14_0, A14B1, n4_14_0);
nor gn6_14_0(n6_14_0, A14B1, n5_14_0);
nor gn7_14_0(n7_14_0, n4_14_0, n5_14_0);
nor gn8_14_0(S14_0, n6_14_0, n7_14_0);
nor gn9_14_0(C14_0, n1_14_0, n5_14_0);

/* FA MFA0_1(S0_1,C0_1,S1_0,C0_0,A0B2); */
nor gn1_0_1(n1_0_1, S1_0, C0_0);
nor gn2_0_1(n2_0_1, n1_0_1, C0_0);
nor gn3_0_1(n3_0_1, S1_0, n1_0_1);
nor gn4_0_1(n4_0_1, n2_0_1, n3_0_1);
nor gn5_0_1(n5_0_1, A0B2, n4_0_1);
nor gn6_0_1(n6_0_1, A0B2, n5_0_1);
nor gn7_0_1(n7_0_1, n4_0_1, n5_0_1);
nor gn8_0_1(S0_1, n6_0_1, n7_0_1);
nor gn9_0_1(C0_1, n1_0_1, n5_0_1);

/* FA MFA1_1(S1_1,C1_1,S2_0,C1_0,A1B2); */
nor gn1_1_1(n1_1_1, S2_0, C1_0);
nor gn2_1_1(n2_1_1, n1_1_1, C1_0);
nor gn3_1_1(n3_1_1, S2_0, n1_1_1);
nor gn4_1_1(n4_1_1, n2_1_1, n3_1_1);
nor gn5_1_1(n5_1_1, A1B2, n4_1_1);
nor gn6_1_1(n6_1_1, A1B2, n5_1_1);
nor gn7_1_1(n7_1_1, n4_1_1, n5_1_1);
nor gn8_1_1(S1_1, n6_1_1, n7_1_1);
nor gn9_1_1(C1_1, n1_1_1, n5_1_1);

/* FA MFA2_1(S2_1,C2_1,S3_0,C2_0,A2B2); */
nor gn1_2_1(n1_2_1, S3_0, C2_0);
nor gn2_2_1(n2_2_1, n1_2_1, C2_0);
nor gn3_2_1(n3_2_1, S3_0, n1_2_1);
nor gn4_2_1(n4_2_1, n2_2_1, n3_2_1);
nor gn5_2_1(n5_2_1, A2B2, n4_2_1);
nor gn6_2_1(n6_2_1, A2B2, n5_2_1);
nor gn7_2_1(n7_2_1, n4_2_1, n5_2_1);
nor gn8_2_1(S2_1, n6_2_1, n7_2_1);
nor gn9_2_1(C2_1, n1_2_1, n5_2_1);

/* FA MFA3_1(S3_1,C3_1,S4_0,C3_0,A3B2); */
nor gn1_3_1(n1_3_1, S4_0, C3_0);
nor gn2_3_1(n2_3_1, n1_3_1, C3_0);
nor gn3_3_1(n3_3_1, S4_0, n1_3_1);
nor gn4_3_1(n4_3_1, n2_3_1, n3_3_1);
nor gn5_3_1(n5_3_1, A3B2, n4_3_1);
nor gn6_3_1(n6_3_1, A3B2, n5_3_1);
nor gn7_3_1(n7_3_1, n4_3_1, n5_3_1);
nor gn8_3_1(S3_1, n6_3_1, n7_3_1);
nor gn9_3_1(C3_1, n1_3_1, n5_3_1);

/* FA MFA4_1(S4_1,C4_1,S5_0,C4_0,A4B2); */
nor gn1_4_1(n1_4_1, S5_0, C4_0);
nor gn2_4_1(n2_4_1, n1_4_1, C4_0);
nor gn3_4_1(n3_4_1, S5_0, n1_4_1);
nor gn4_4_1(n4_4_1, n2_4_1, n3_4_1);
nor gn5_4_1(n5_4_1, A4B2, n4_4_1);
nor gn6_4_1(n6_4_1, A4B2, n5_4_1);
nor gn7_4_1(n7_4_1, n4_4_1, n5_4_1);
nor gn8_4_1(S4_1, n6_4_1, n7_4_1);
nor gn9_4_1(C4_1, n1_4_1, n5_4_1);

/* FA MFA5_1(S5_1,C5_1,S6_0,C5_0,A5B2); */
nor gn1_5_1(n1_5_1, S6_0, C5_0);
nor gn2_5_1(n2_5_1, n1_5_1, C5_0);
nor gn3_5_1(n3_5_1, S6_0, n1_5_1);
nor gn4_5_1(n4_5_1, n2_5_1, n3_5_1);
nor gn5_5_1(n5_5_1, A5B2, n4_5_1);
nor gn6_5_1(n6_5_1, A5B2, n5_5_1);
nor gn7_5_1(n7_5_1, n4_5_1, n5_5_1);
nor gn8_5_1(S5_1, n6_5_1, n7_5_1);
nor gn9_5_1(C5_1, n1_5_1, n5_5_1);

/* FA MFA6_1(S6_1,C6_1,S7_0,C6_0,A6B2); */
nor gn1_6_1(n1_6_1, S7_0, C6_0);
nor gn2_6_1(n2_6_1, n1_6_1, C6_0);
nor gn3_6_1(n3_6_1, S7_0, n1_6_1);
nor gn4_6_1(n4_6_1, n2_6_1, n3_6_1);
nor gn5_6_1(n5_6_1, A6B2, n4_6_1);
nor gn6_6_1(n6_6_1, A6B2, n5_6_1);
nor gn7_6_1(n7_6_1, n4_6_1, n5_6_1);
nor gn8_6_1(S6_1, n6_6_1, n7_6_1);
nor gn9_6_1(C6_1, n1_6_1, n5_6_1);

/* FA MFA7_1(S7_1,C7_1,S8_0,C7_0,A7B2); */
nor gn1_7_1(n1_7_1, S8_0, C7_0);
nor gn2_7_1(n2_7_1, n1_7_1, C7_0);
nor gn3_7_1(n3_7_1, S8_0, n1_7_1);
nor gn4_7_1(n4_7_1, n2_7_1, n3_7_1);
nor gn5_7_1(n5_7_1, A7B2, n4_7_1);
nor gn6_7_1(n6_7_1, A7B2, n5_7_1);
nor gn7_7_1(n7_7_1, n4_7_1, n5_7_1);
nor gn8_7_1(S7_1, n6_7_1, n7_7_1);
nor gn9_7_1(C7_1, n1_7_1, n5_7_1);

/* FA MFA8_1(S8_1,C8_1,S9_0,C8_0,A8B2); */
nor gn1_8_1(n1_8_1, S9_0, C8_0);
nor gn2_8_1(n2_8_1, n1_8_1, C8_0);
nor gn3_8_1(n3_8_1, S9_0, n1_8_1);
nor gn4_8_1(n4_8_1, n2_8_1, n3_8_1);
nor gn5_8_1(n5_8_1, A8B2, n4_8_1);
nor gn6_8_1(n6_8_1, A8B2, n5_8_1);
nor gn7_8_1(n7_8_1, n4_8_1, n5_8_1);
nor gn8_8_1(S8_1, n6_8_1, n7_8_1);
nor gn9_8_1(C8_1, n1_8_1, n5_8_1);

/* FA MFA9_1(S9_1,C9_1,S10_0,C9_0,A9B2); */
nor gn1_9_1(n1_9_1, S10_0, C9_0);
nor gn2_9_1(n2_9_1, n1_9_1, C9_0);
nor gn3_9_1(n3_9_1, S10_0, n1_9_1);
nor gn4_9_1(n4_9_1, n2_9_1, n3_9_1);
nor gn5_9_1(n5_9_1, A9B2, n4_9_1);
nor gn6_9_1(n6_9_1, A9B2, n5_9_1);
nor gn7_9_1(n7_9_1, n4_9_1, n5_9_1);
nor gn8_9_1(S9_1, n6_9_1, n7_9_1);
nor gn9_9_1(C9_1, n1_9_1, n5_9_1);

/* FA MFA10_1(S10_1,C10_1,S11_0,C10_0,A10B2); */
nor gn1_10_1(n1_10_1, S11_0, C10_0);
nor gn2_10_1(n2_10_1, n1_10_1, C10_0);
nor gn3_10_1(n3_10_1, S11_0, n1_10_1);
nor gn4_10_1(n4_10_1, n2_10_1, n3_10_1);
nor gn5_10_1(n5_10_1, A10B2, n4_10_1);
nor gn6_10_1(n6_10_1, A10B2, n5_10_1);
nor gn7_10_1(n7_10_1, n4_10_1, n5_10_1);
nor gn8_10_1(S10_1, n6_10_1, n7_10_1);
nor gn9_10_1(C10_1, n1_10_1, n5_10_1);

/* FA MFA11_1(S11_1,C11_1,S12_0,C11_0,A11B2); */
nor gn1_11_1(n1_11_1, S12_0, C11_0);
nor gn2_11_1(n2_11_1, n1_11_1, C11_0);
nor gn3_11_1(n3_11_1, S12_0, n1_11_1);
nor gn4_11_1(n4_11_1, n2_11_1, n3_11_1);
nor gn5_11_1(n5_11_1, A11B2, n4_11_1);
nor gn6_11_1(n6_11_1, A11B2, n5_11_1);
nor gn7_11_1(n7_11_1, n4_11_1, n5_11_1);
nor gn8_11_1(S11_1, n6_11_1, n7_11_1);
nor gn9_11_1(C11_1, n1_11_1, n5_11_1);

/* FA MFA12_1(S12_1,C12_1,S13_0,C12_0,A12B2); */
nor gn1_12_1(n1_12_1, S13_0, C12_0);
nor gn2_12_1(n2_12_1, n1_12_1, C12_0);
nor gn3_12_1(n3_12_1, S13_0, n1_12_1);
nor gn4_12_1(n4_12_1, n2_12_1, n3_12_1);
nor gn5_12_1(n5_12_1, A12B2, n4_12_1);
nor gn6_12_1(n6_12_1, A12B2, n5_12_1);
nor gn7_12_1(n7_12_1, n4_12_1, n5_12_1);
nor gn8_12_1(S12_1, n6_12_1, n7_12_1);
nor gn9_12_1(C12_1, n1_12_1, n5_12_1);

/* FA MFA13_1(S13_1,C13_1,S14_0,C13_0,A13B2); */
nor gn1_13_1(n1_13_1, S14_0, C13_0);
nor gn2_13_1(n2_13_1, n1_13_1, C13_0);
nor gn3_13_1(n3_13_1, S14_0, n1_13_1);
nor gn4_13_1(n4_13_1, n2_13_1, n3_13_1);
nor gn5_13_1(n5_13_1, A13B2, n4_13_1);
nor gn6_13_1(n6_13_1, A13B2, n5_13_1);
nor gn7_13_1(n7_13_1, n4_13_1, n5_13_1);
nor gn8_13_1(S13_1, n6_13_1, n7_13_1);
nor gn9_13_1(C13_1, n1_13_1, n5_13_1);

/* FA MFA14_1(S14_1,C14_1,A15B1,C14_0,A14B2); */
nor gn1_14_1(n1_14_1, A15B1, C14_0);
nor gn2_14_1(n2_14_1, n1_14_1, C14_0);
nor gn3_14_1(n3_14_1, A15B1, n1_14_1);
nor gn4_14_1(n4_14_1, n2_14_1, n3_14_1);
nor gn5_14_1(n5_14_1, A14B2, n4_14_1);
nor gn6_14_1(n6_14_1, A14B2, n5_14_1);
nor gn7_14_1(n7_14_1, n4_14_1, n5_14_1);
nor gn8_14_1(S14_1, n6_14_1, n7_14_1);
nor gn9_14_1(C14_1, n1_14_1, n5_14_1);

/* FA MFA0_2(S0_2,C0_2,S1_1,C0_1,A0B3); */
nor gn1_0_2(n1_0_2, S1_1, C0_1);
nor gn2_0_2(n2_0_2, n1_0_2, C0_1);
nor gn3_0_2(n3_0_2, S1_1, n1_0_2);
nor gn4_0_2(n4_0_2, n2_0_2, n3_0_2);
nor gn5_0_2(n5_0_2, A0B3, n4_0_2);
nor gn6_0_2(n6_0_2, A0B3, n5_0_2);
nor gn7_0_2(n7_0_2, n4_0_2, n5_0_2);
nor gn8_0_2(S0_2, n6_0_2, n7_0_2);
nor gn9_0_2(C0_2, n1_0_2, n5_0_2);

/* FA MFA1_2(S1_2,C1_2,S2_1,C1_1,A1B3); */
nor gn1_1_2(n1_1_2, S2_1, C1_1);
nor gn2_1_2(n2_1_2, n1_1_2, C1_1);
nor gn3_1_2(n3_1_2, S2_1, n1_1_2);
nor gn4_1_2(n4_1_2, n2_1_2, n3_1_2);
nor gn5_1_2(n5_1_2, A1B3, n4_1_2);
nor gn6_1_2(n6_1_2, A1B3, n5_1_2);
nor gn7_1_2(n7_1_2, n4_1_2, n5_1_2);
nor gn8_1_2(S1_2, n6_1_2, n7_1_2);
nor gn9_1_2(C1_2, n1_1_2, n5_1_2);

/* FA MFA2_2(S2_2,C2_2,S3_1,C2_1,A2B3); */
nor gn1_2_2(n1_2_2, S3_1, C2_1);
nor gn2_2_2(n2_2_2, n1_2_2, C2_1);
nor gn3_2_2(n3_2_2, S3_1, n1_2_2);
nor gn4_2_2(n4_2_2, n2_2_2, n3_2_2);
nor gn5_2_2(n5_2_2, A2B3, n4_2_2);
nor gn6_2_2(n6_2_2, A2B3, n5_2_2);
nor gn7_2_2(n7_2_2, n4_2_2, n5_2_2);
nor gn8_2_2(S2_2, n6_2_2, n7_2_2);
nor gn9_2_2(C2_2, n1_2_2, n5_2_2);

/* FA MFA3_2(S3_2,C3_2,S4_1,C3_1,A3B3); */
nor gn1_3_2(n1_3_2, S4_1, C3_1);
nor gn2_3_2(n2_3_2, n1_3_2, C3_1);
nor gn3_3_2(n3_3_2, S4_1, n1_3_2);
nor gn4_3_2(n4_3_2, n2_3_2, n3_3_2);
nor gn5_3_2(n5_3_2, A3B3, n4_3_2);
nor gn6_3_2(n6_3_2, A3B3, n5_3_2);
nor gn7_3_2(n7_3_2, n4_3_2, n5_3_2);
nor gn8_3_2(S3_2, n6_3_2, n7_3_2);
nor gn9_3_2(C3_2, n1_3_2, n5_3_2);

/* FA MFA4_2(S4_2,C4_2,S5_1,C4_1,A4B3); */
nor gn1_4_2(n1_4_2, S5_1, C4_1);
nor gn2_4_2(n2_4_2, n1_4_2, C4_1);
nor gn3_4_2(n3_4_2, S5_1, n1_4_2);
nor gn4_4_2(n4_4_2, n2_4_2, n3_4_2);
nor gn5_4_2(n5_4_2, A4B3, n4_4_2);
nor gn6_4_2(n6_4_2, A4B3, n5_4_2);
nor gn7_4_2(n7_4_2, n4_4_2, n5_4_2);
nor gn8_4_2(S4_2, n6_4_2, n7_4_2);
nor gn9_4_2(C4_2, n1_4_2, n5_4_2);

/* FA MFA5_2(S5_2,C5_2,S6_1,C5_1,A5B3); */
nor gn1_5_2(n1_5_2, S6_1, C5_1);
nor gn2_5_2(n2_5_2, n1_5_2, C5_1);
nor gn3_5_2(n3_5_2, S6_1, n1_5_2);
nor gn4_5_2(n4_5_2, n2_5_2, n3_5_2);
nor gn5_5_2(n5_5_2, A5B3, n4_5_2);
nor gn6_5_2(n6_5_2, A5B3, n5_5_2);
nor gn7_5_2(n7_5_2, n4_5_2, n5_5_2);
nor gn8_5_2(S5_2, n6_5_2, n7_5_2);
nor gn9_5_2(C5_2, n1_5_2, n5_5_2);

/* FA MFA6_2(S6_2,C6_2,S7_1,C6_1,A6B3); */
nor gn1_6_2(n1_6_2, S7_1, C6_1);
nor gn2_6_2(n2_6_2, n1_6_2, C6_1);
nor gn3_6_2(n3_6_2, S7_1, n1_6_2);
nor gn4_6_2(n4_6_2, n2_6_2, n3_6_2);
nor gn5_6_2(n5_6_2, A6B3, n4_6_2);
nor gn6_6_2(n6_6_2, A6B3, n5_6_2);
nor gn7_6_2(n7_6_2, n4_6_2, n5_6_2);
nor gn8_6_2(S6_2, n6_6_2, n7_6_2);
nor gn9_6_2(C6_2, n1_6_2, n5_6_2);

/* FA MFA7_2(S7_2,C7_2,S8_1,C7_1,A7B3); */
nor gn1_7_2(n1_7_2, S8_1, C7_1);
nor gn2_7_2(n2_7_2, n1_7_2, C7_1);
nor gn3_7_2(n3_7_2, S8_1, n1_7_2);
nor gn4_7_2(n4_7_2, n2_7_2, n3_7_2);
nor gn5_7_2(n5_7_2, A7B3, n4_7_2);
nor gn6_7_2(n6_7_2, A7B3, n5_7_2);
nor gn7_7_2(n7_7_2, n4_7_2, n5_7_2);
nor gn8_7_2(S7_2, n6_7_2, n7_7_2);
nor gn9_7_2(C7_2, n1_7_2, n5_7_2);

/* FA MFA8_2(S8_2,C8_2,S9_1,C8_1,A8B3); */
nor gn1_8_2(n1_8_2, S9_1, C8_1);
nor gn2_8_2(n2_8_2, n1_8_2, C8_1);
nor gn3_8_2(n3_8_2, S9_1, n1_8_2);
nor gn4_8_2(n4_8_2, n2_8_2, n3_8_2);
nor gn5_8_2(n5_8_2, A8B3, n4_8_2);
nor gn6_8_2(n6_8_2, A8B3, n5_8_2);
nor gn7_8_2(n7_8_2, n4_8_2, n5_8_2);
nor gn8_8_2(S8_2, n6_8_2, n7_8_2);
nor gn9_8_2(C8_2, n1_8_2, n5_8_2);

/* FA MFA9_2(S9_2,C9_2,S10_1,C9_1,A9B3); */
nor gn1_9_2(n1_9_2, S10_1, C9_1);
nor gn2_9_2(n2_9_2, n1_9_2, C9_1);
nor gn3_9_2(n3_9_2, S10_1, n1_9_2);
nor gn4_9_2(n4_9_2, n2_9_2, n3_9_2);
nor gn5_9_2(n5_9_2, A9B3, n4_9_2);
nor gn6_9_2(n6_9_2, A9B3, n5_9_2);
nor gn7_9_2(n7_9_2, n4_9_2, n5_9_2);
nor gn8_9_2(S9_2, n6_9_2, n7_9_2);
nor gn9_9_2(C9_2, n1_9_2, n5_9_2);

/* FA MFA10_2(S10_2,C10_2,S11_1,C10_1,A10B3); */
nor gn1_10_2(n1_10_2, S11_1, C10_1);
nor gn2_10_2(n2_10_2, n1_10_2, C10_1);
nor gn3_10_2(n3_10_2, S11_1, n1_10_2);
nor gn4_10_2(n4_10_2, n2_10_2, n3_10_2);
nor gn5_10_2(n5_10_2, A10B3, n4_10_2);
nor gn6_10_2(n6_10_2, A10B3, n5_10_2);
nor gn7_10_2(n7_10_2, n4_10_2, n5_10_2);
nor gn8_10_2(S10_2, n6_10_2, n7_10_2);
nor gn9_10_2(C10_2, n1_10_2, n5_10_2);

/* FA MFA11_2(S11_2,C11_2,S12_1,C11_1,A11B3); */
nor gn1_11_2(n1_11_2, S12_1, C11_1);
nor gn2_11_2(n2_11_2, n1_11_2, C11_1);
nor gn3_11_2(n3_11_2, S12_1, n1_11_2);
nor gn4_11_2(n4_11_2, n2_11_2, n3_11_2);
nor gn5_11_2(n5_11_2, A11B3, n4_11_2);
nor gn6_11_2(n6_11_2, A11B3, n5_11_2);
nor gn7_11_2(n7_11_2, n4_11_2, n5_11_2);
nor gn8_11_2(S11_2, n6_11_2, n7_11_2);
nor gn9_11_2(C11_2, n1_11_2, n5_11_2);

/* FA MFA12_2(S12_2,C12_2,S13_1,C12_1,A12B3); */
nor gn1_12_2(n1_12_2, S13_1, C12_1);
nor gn2_12_2(n2_12_2, n1_12_2, C12_1);
nor gn3_12_2(n3_12_2, S13_1, n1_12_2);
nor gn4_12_2(n4_12_2, n2_12_2, n3_12_2);
nor gn5_12_2(n5_12_2, A12B3, n4_12_2);
nor gn6_12_2(n6_12_2, A12B3, n5_12_2);
nor gn7_12_2(n7_12_2, n4_12_2, n5_12_2);
nor gn8_12_2(S12_2, n6_12_2, n7_12_2);
nor gn9_12_2(C12_2, n1_12_2, n5_12_2);

/* FA MFA13_2(S13_2,C13_2,S14_1,C13_1,A13B3); */
nor gn1_13_2(n1_13_2, S14_1, C13_1);
nor gn2_13_2(n2_13_2, n1_13_2, C13_1);
nor gn3_13_2(n3_13_2, S14_1, n1_13_2);
nor gn4_13_2(n4_13_2, n2_13_2, n3_13_2);
nor gn5_13_2(n5_13_2, A13B3, n4_13_2);
nor gn6_13_2(n6_13_2, A13B3, n5_13_2);
nor gn7_13_2(n7_13_2, n4_13_2, n5_13_2);
nor gn8_13_2(S13_2, n6_13_2, n7_13_2);
nor gn9_13_2(C13_2, n1_13_2, n5_13_2);

/* FA MFA14_2(S14_2,C14_2,A15B2,C14_1,A14B3); */
nor gn1_14_2(n1_14_2, A15B2, C14_1);
nor gn2_14_2(n2_14_2, n1_14_2, C14_1);
nor gn3_14_2(n3_14_2, A15B2, n1_14_2);
nor gn4_14_2(n4_14_2, n2_14_2, n3_14_2);
nor gn5_14_2(n5_14_2, A14B3, n4_14_2);
nor gn6_14_2(n6_14_2, A14B3, n5_14_2);
nor gn7_14_2(n7_14_2, n4_14_2, n5_14_2);
nor gn8_14_2(S14_2, n6_14_2, n7_14_2);
nor gn9_14_2(C14_2, n1_14_2, n5_14_2);

/* FA MFA0_3(S0_3,C0_3,S1_2,C0_2,A0B4); */
nor gn1_0_3(n1_0_3, S1_2, C0_2);
nor gn2_0_3(n2_0_3, n1_0_3, C0_2);
nor gn3_0_3(n3_0_3, S1_2, n1_0_3);
nor gn4_0_3(n4_0_3, n2_0_3, n3_0_3);
nor gn5_0_3(n5_0_3, A0B4, n4_0_3);
nor gn6_0_3(n6_0_3, A0B4, n5_0_3);
nor gn7_0_3(n7_0_3, n4_0_3, n5_0_3);
nor gn8_0_3(S0_3, n6_0_3, n7_0_3);
nor gn9_0_3(C0_3, n1_0_3, n5_0_3);

/* FA MFA1_3(S1_3,C1_3,S2_2,C1_2,A1B4); */
nor gn1_1_3(n1_1_3, S2_2, C1_2);
nor gn2_1_3(n2_1_3, n1_1_3, C1_2);
nor gn3_1_3(n3_1_3, S2_2, n1_1_3);
nor gn4_1_3(n4_1_3, n2_1_3, n3_1_3);
nor gn5_1_3(n5_1_3, A1B4, n4_1_3);
nor gn6_1_3(n6_1_3, A1B4, n5_1_3);
nor gn7_1_3(n7_1_3, n4_1_3, n5_1_3);
nor gn8_1_3(S1_3, n6_1_3, n7_1_3);
nor gn9_1_3(C1_3, n1_1_3, n5_1_3);

/* FA MFA2_3(S2_3,C2_3,S3_2,C2_2,A2B4); */
nor gn1_2_3(n1_2_3, S3_2, C2_2);
nor gn2_2_3(n2_2_3, n1_2_3, C2_2);
nor gn3_2_3(n3_2_3, S3_2, n1_2_3);
nor gn4_2_3(n4_2_3, n2_2_3, n3_2_3);
nor gn5_2_3(n5_2_3, A2B4, n4_2_3);
nor gn6_2_3(n6_2_3, A2B4, n5_2_3);
nor gn7_2_3(n7_2_3, n4_2_3, n5_2_3);
nor gn8_2_3(S2_3, n6_2_3, n7_2_3);
nor gn9_2_3(C2_3, n1_2_3, n5_2_3);

/* FA MFA3_3(S3_3,C3_3,S4_2,C3_2,A3B4); */
nor gn1_3_3(n1_3_3, S4_2, C3_2);
nor gn2_3_3(n2_3_3, n1_3_3, C3_2);
nor gn3_3_3(n3_3_3, S4_2, n1_3_3);
nor gn4_3_3(n4_3_3, n2_3_3, n3_3_3);
nor gn5_3_3(n5_3_3, A3B4, n4_3_3);
nor gn6_3_3(n6_3_3, A3B4, n5_3_3);
nor gn7_3_3(n7_3_3, n4_3_3, n5_3_3);
nor gn8_3_3(S3_3, n6_3_3, n7_3_3);
nor gn9_3_3(C3_3, n1_3_3, n5_3_3);

/* FA MFA4_3(S4_3,C4_3,S5_2,C4_2,A4B4); */
nor gn1_4_3(n1_4_3, S5_2, C4_2);
nor gn2_4_3(n2_4_3, n1_4_3, C4_2);
nor gn3_4_3(n3_4_3, S5_2, n1_4_3);
nor gn4_4_3(n4_4_3, n2_4_3, n3_4_3);
nor gn5_4_3(n5_4_3, A4B4, n4_4_3);
nor gn6_4_3(n6_4_3, A4B4, n5_4_3);
nor gn7_4_3(n7_4_3, n4_4_3, n5_4_3);
nor gn8_4_3(S4_3, n6_4_3, n7_4_3);
nor gn9_4_3(C4_3, n1_4_3, n5_4_3);

/* FA MFA5_3(S5_3,C5_3,S6_2,C5_2,A5B4); */
nor gn1_5_3(n1_5_3, S6_2, C5_2);
nor gn2_5_3(n2_5_3, n1_5_3, C5_2);
nor gn3_5_3(n3_5_3, S6_2, n1_5_3);
nor gn4_5_3(n4_5_3, n2_5_3, n3_5_3);
nor gn5_5_3(n5_5_3, A5B4, n4_5_3);
nor gn6_5_3(n6_5_3, A5B4, n5_5_3);
nor gn7_5_3(n7_5_3, n4_5_3, n5_5_3);
nor gn8_5_3(S5_3, n6_5_3, n7_5_3);
nor gn9_5_3(C5_3, n1_5_3, n5_5_3);

/* FA MFA6_3(S6_3,C6_3,S7_2,C6_2,A6B4); */
nor gn1_6_3(n1_6_3, S7_2, C6_2);
nor gn2_6_3(n2_6_3, n1_6_3, C6_2);
nor gn3_6_3(n3_6_3, S7_2, n1_6_3);
nor gn4_6_3(n4_6_3, n2_6_3, n3_6_3);
nor gn5_6_3(n5_6_3, A6B4, n4_6_3);
nor gn6_6_3(n6_6_3, A6B4, n5_6_3);
nor gn7_6_3(n7_6_3, n4_6_3, n5_6_3);
nor gn8_6_3(S6_3, n6_6_3, n7_6_3);
nor gn9_6_3(C6_3, n1_6_3, n5_6_3);

/* FA MFA7_3(S7_3,C7_3,S8_2,C7_2,A7B4); */
nor gn1_7_3(n1_7_3, S8_2, C7_2);
nor gn2_7_3(n2_7_3, n1_7_3, C7_2);
nor gn3_7_3(n3_7_3, S8_2, n1_7_3);
nor gn4_7_3(n4_7_3, n2_7_3, n3_7_3);
nor gn5_7_3(n5_7_3, A7B4, n4_7_3);
nor gn6_7_3(n6_7_3, A7B4, n5_7_3);
nor gn7_7_3(n7_7_3, n4_7_3, n5_7_3);
nor gn8_7_3(S7_3, n6_7_3, n7_7_3);
nor gn9_7_3(C7_3, n1_7_3, n5_7_3);

/* FA MFA8_3(S8_3,C8_3,S9_2,C8_2,A8B4); */
nor gn1_8_3(n1_8_3, S9_2, C8_2);
nor gn2_8_3(n2_8_3, n1_8_3, C8_2);
nor gn3_8_3(n3_8_3, S9_2, n1_8_3);
nor gn4_8_3(n4_8_3, n2_8_3, n3_8_3);
nor gn5_8_3(n5_8_3, A8B4, n4_8_3);
nor gn6_8_3(n6_8_3, A8B4, n5_8_3);
nor gn7_8_3(n7_8_3, n4_8_3, n5_8_3);
nor gn8_8_3(S8_3, n6_8_3, n7_8_3);
nor gn9_8_3(C8_3, n1_8_3, n5_8_3);

/* FA MFA9_3(S9_3,C9_3,S10_2,C9_2,A9B4); */
nor gn1_9_3(n1_9_3, S10_2, C9_2);
nor gn2_9_3(n2_9_3, n1_9_3, C9_2);
nor gn3_9_3(n3_9_3, S10_2, n1_9_3);
nor gn4_9_3(n4_9_3, n2_9_3, n3_9_3);
nor gn5_9_3(n5_9_3, A9B4, n4_9_3);
nor gn6_9_3(n6_9_3, A9B4, n5_9_3);
nor gn7_9_3(n7_9_3, n4_9_3, n5_9_3);
nor gn8_9_3(S9_3, n6_9_3, n7_9_3);
nor gn9_9_3(C9_3, n1_9_3, n5_9_3);

/* FA MFA10_3(S10_3,C10_3,S11_2,C10_2,A10B4); */
nor gn1_10_3(n1_10_3, S11_2, C10_2);
nor gn2_10_3(n2_10_3, n1_10_3, C10_2);
nor gn3_10_3(n3_10_3, S11_2, n1_10_3);
nor gn4_10_3(n4_10_3, n2_10_3, n3_10_3);
nor gn5_10_3(n5_10_3, A10B4, n4_10_3);
nor gn6_10_3(n6_10_3, A10B4, n5_10_3);
nor gn7_10_3(n7_10_3, n4_10_3, n5_10_3);
nor gn8_10_3(S10_3, n6_10_3, n7_10_3);
nor gn9_10_3(C10_3, n1_10_3, n5_10_3);

/* FA MFA11_3(S11_3,C11_3,S12_2,C11_2,A11B4); */
nor gn1_11_3(n1_11_3, S12_2, C11_2);
nor gn2_11_3(n2_11_3, n1_11_3, C11_2);
nor gn3_11_3(n3_11_3, S12_2, n1_11_3);
nor gn4_11_3(n4_11_3, n2_11_3, n3_11_3);
nor gn5_11_3(n5_11_3, A11B4, n4_11_3);
nor gn6_11_3(n6_11_3, A11B4, n5_11_3);
nor gn7_11_3(n7_11_3, n4_11_3, n5_11_3);
nor gn8_11_3(S11_3, n6_11_3, n7_11_3);
nor gn9_11_3(C11_3, n1_11_3, n5_11_3);

/* FA MFA12_3(S12_3,C12_3,S13_2,C12_2,A12B4); */
nor gn1_12_3(n1_12_3, S13_2, C12_2);
nor gn2_12_3(n2_12_3, n1_12_3, C12_2);
nor gn3_12_3(n3_12_3, S13_2, n1_12_3);
nor gn4_12_3(n4_12_3, n2_12_3, n3_12_3);
nor gn5_12_3(n5_12_3, A12B4, n4_12_3);
nor gn6_12_3(n6_12_3, A12B4, n5_12_3);
nor gn7_12_3(n7_12_3, n4_12_3, n5_12_3);
nor gn8_12_3(S12_3, n6_12_3, n7_12_3);
nor gn9_12_3(C12_3, n1_12_3, n5_12_3);

/* FA MFA13_3(S13_3,C13_3,S14_2,C13_2,A13B4); */
nor gn1_13_3(n1_13_3, S14_2, C13_2);
nor gn2_13_3(n2_13_3, n1_13_3, C13_2);
nor gn3_13_3(n3_13_3, S14_2, n1_13_3);
nor gn4_13_3(n4_13_3, n2_13_3, n3_13_3);
nor gn5_13_3(n5_13_3, A13B4, n4_13_3);
nor gn6_13_3(n6_13_3, A13B4, n5_13_3);
nor gn7_13_3(n7_13_3, n4_13_3, n5_13_3);
nor gn8_13_3(S13_3, n6_13_3, n7_13_3);
nor gn9_13_3(C13_3, n1_13_3, n5_13_3);

/* FA MFA14_3(S14_3,C14_3,A15B3,C14_2,A14B4); */
nor gn1_14_3(n1_14_3, A15B3, C14_2);
nor gn2_14_3(n2_14_3, n1_14_3, C14_2);
nor gn3_14_3(n3_14_3, A15B3, n1_14_3);
nor gn4_14_3(n4_14_3, n2_14_3, n3_14_3);
nor gn5_14_3(n5_14_3, A14B4, n4_14_3);
nor gn6_14_3(n6_14_3, A14B4, n5_14_3);
nor gn7_14_3(n7_14_3, n4_14_3, n5_14_3);
nor gn8_14_3(S14_3, n6_14_3, n7_14_3);
nor gn9_14_3(C14_3, n1_14_3, n5_14_3);

/* FA MFA0_4(S0_4,C0_4,S1_3,C0_3,A0B5); */
nor gn1_0_4(n1_0_4, S1_3, C0_3);
nor gn2_0_4(n2_0_4, n1_0_4, C0_3);
nor gn3_0_4(n3_0_4, S1_3, n1_0_4);
nor gn4_0_4(n4_0_4, n2_0_4, n3_0_4);
nor gn5_0_4(n5_0_4, A0B5, n4_0_4);
nor gn6_0_4(n6_0_4, A0B5, n5_0_4);
nor gn7_0_4(n7_0_4, n4_0_4, n5_0_4);
nor gn8_0_4(S0_4, n6_0_4, n7_0_4);
nor gn9_0_4(C0_4, n1_0_4, n5_0_4);

/* FA MFA1_4(S1_4,C1_4,S2_3,C1_3,A1B5); */
nor gn1_1_4(n1_1_4, S2_3, C1_3);
nor gn2_1_4(n2_1_4, n1_1_4, C1_3);
nor gn3_1_4(n3_1_4, S2_3, n1_1_4);
nor gn4_1_4(n4_1_4, n2_1_4, n3_1_4);
nor gn5_1_4(n5_1_4, A1B5, n4_1_4);
nor gn6_1_4(n6_1_4, A1B5, n5_1_4);
nor gn7_1_4(n7_1_4, n4_1_4, n5_1_4);
nor gn8_1_4(S1_4, n6_1_4, n7_1_4);
nor gn9_1_4(C1_4, n1_1_4, n5_1_4);

/* FA MFA2_4(S2_4,C2_4,S3_3,C2_3,A2B5); */
nor gn1_2_4(n1_2_4, S3_3, C2_3);
nor gn2_2_4(n2_2_4, n1_2_4, C2_3);
nor gn3_2_4(n3_2_4, S3_3, n1_2_4);
nor gn4_2_4(n4_2_4, n2_2_4, n3_2_4);
nor gn5_2_4(n5_2_4, A2B5, n4_2_4);
nor gn6_2_4(n6_2_4, A2B5, n5_2_4);
nor gn7_2_4(n7_2_4, n4_2_4, n5_2_4);
nor gn8_2_4(S2_4, n6_2_4, n7_2_4);
nor gn9_2_4(C2_4, n1_2_4, n5_2_4);

/* FA MFA3_4(S3_4,C3_4,S4_3,C3_3,A3B5); */
nor gn1_3_4(n1_3_4, S4_3, C3_3);
nor gn2_3_4(n2_3_4, n1_3_4, C3_3);
nor gn3_3_4(n3_3_4, S4_3, n1_3_4);
nor gn4_3_4(n4_3_4, n2_3_4, n3_3_4);
nor gn5_3_4(n5_3_4, A3B5, n4_3_4);
nor gn6_3_4(n6_3_4, A3B5, n5_3_4);
nor gn7_3_4(n7_3_4, n4_3_4, n5_3_4);
nor gn8_3_4(S3_4, n6_3_4, n7_3_4);
nor gn9_3_4(C3_4, n1_3_4, n5_3_4);

/* FA MFA4_4(S4_4,C4_4,S5_3,C4_3,A4B5); */
nor gn1_4_4(n1_4_4, S5_3, C4_3);
nor gn2_4_4(n2_4_4, n1_4_4, C4_3);
nor gn3_4_4(n3_4_4, S5_3, n1_4_4);
nor gn4_4_4(n4_4_4, n2_4_4, n3_4_4);
nor gn5_4_4(n5_4_4, A4B5, n4_4_4);
nor gn6_4_4(n6_4_4, A4B5, n5_4_4);
nor gn7_4_4(n7_4_4, n4_4_4, n5_4_4);
nor gn8_4_4(S4_4, n6_4_4, n7_4_4);
nor gn9_4_4(C4_4, n1_4_4, n5_4_4);

/* FA MFA5_4(S5_4,C5_4,S6_3,C5_3,A5B5); */
nor gn1_5_4(n1_5_4, S6_3, C5_3);
nor gn2_5_4(n2_5_4, n1_5_4, C5_3);
nor gn3_5_4(n3_5_4, S6_3, n1_5_4);
nor gn4_5_4(n4_5_4, n2_5_4, n3_5_4);
nor gn5_5_4(n5_5_4, A5B5, n4_5_4);
nor gn6_5_4(n6_5_4, A5B5, n5_5_4);
nor gn7_5_4(n7_5_4, n4_5_4, n5_5_4);
nor gn8_5_4(S5_4, n6_5_4, n7_5_4);
nor gn9_5_4(C5_4, n1_5_4, n5_5_4);

/* FA MFA6_4(S6_4,C6_4,S7_3,C6_3,A6B5); */
nor gn1_6_4(n1_6_4, S7_3, C6_3);
nor gn2_6_4(n2_6_4, n1_6_4, C6_3);
nor gn3_6_4(n3_6_4, S7_3, n1_6_4);
nor gn4_6_4(n4_6_4, n2_6_4, n3_6_4);
nor gn5_6_4(n5_6_4, A6B5, n4_6_4);
nor gn6_6_4(n6_6_4, A6B5, n5_6_4);
nor gn7_6_4(n7_6_4, n4_6_4, n5_6_4);
nor gn8_6_4(S6_4, n6_6_4, n7_6_4);
nor gn9_6_4(C6_4, n1_6_4, n5_6_4);

/* FA MFA7_4(S7_4,C7_4,S8_3,C7_3,A7B5); */
nor gn1_7_4(n1_7_4, S8_3, C7_3);
nor gn2_7_4(n2_7_4, n1_7_4, C7_3);
nor gn3_7_4(n3_7_4, S8_3, n1_7_4);
nor gn4_7_4(n4_7_4, n2_7_4, n3_7_4);
nor gn5_7_4(n5_7_4, A7B5, n4_7_4);
nor gn6_7_4(n6_7_4, A7B5, n5_7_4);
nor gn7_7_4(n7_7_4, n4_7_4, n5_7_4);
nor gn8_7_4(S7_4, n6_7_4, n7_7_4);
nor gn9_7_4(C7_4, n1_7_4, n5_7_4);

/* FA MFA8_4(S8_4,C8_4,S9_3,C8_3,A8B5); */
nor gn1_8_4(n1_8_4, S9_3, C8_3);
nor gn2_8_4(n2_8_4, n1_8_4, C8_3);
nor gn3_8_4(n3_8_4, S9_3, n1_8_4);
nor gn4_8_4(n4_8_4, n2_8_4, n3_8_4);
nor gn5_8_4(n5_8_4, A8B5, n4_8_4);
nor gn6_8_4(n6_8_4, A8B5, n5_8_4);
nor gn7_8_4(n7_8_4, n4_8_4, n5_8_4);
nor gn8_8_4(S8_4, n6_8_4, n7_8_4);
nor gn9_8_4(C8_4, n1_8_4, n5_8_4);

/* FA MFA9_4(S9_4,C9_4,S10_3,C9_3,A9B5); */
nor gn1_9_4(n1_9_4, S10_3, C9_3);
nor gn2_9_4(n2_9_4, n1_9_4, C9_3);
nor gn3_9_4(n3_9_4, S10_3, n1_9_4);
nor gn4_9_4(n4_9_4, n2_9_4, n3_9_4);
nor gn5_9_4(n5_9_4, A9B5, n4_9_4);
nor gn6_9_4(n6_9_4, A9B5, n5_9_4);
nor gn7_9_4(n7_9_4, n4_9_4, n5_9_4);
nor gn8_9_4(S9_4, n6_9_4, n7_9_4);
nor gn9_9_4(C9_4, n1_9_4, n5_9_4);

/* FA MFA10_4(S10_4,C10_4,S11_3,C10_3,A10B5); */
nor gn1_10_4(n1_10_4, S11_3, C10_3);
nor gn2_10_4(n2_10_4, n1_10_4, C10_3);
nor gn3_10_4(n3_10_4, S11_3, n1_10_4);
nor gn4_10_4(n4_10_4, n2_10_4, n3_10_4);
nor gn5_10_4(n5_10_4, A10B5, n4_10_4);
nor gn6_10_4(n6_10_4, A10B5, n5_10_4);
nor gn7_10_4(n7_10_4, n4_10_4, n5_10_4);
nor gn8_10_4(S10_4, n6_10_4, n7_10_4);
nor gn9_10_4(C10_4, n1_10_4, n5_10_4);

/* FA MFA11_4(S11_4,C11_4,S12_3,C11_3,A11B5); */
nor gn1_11_4(n1_11_4, S12_3, C11_3);
nor gn2_11_4(n2_11_4, n1_11_4, C11_3);
nor gn3_11_4(n3_11_4, S12_3, n1_11_4);
nor gn4_11_4(n4_11_4, n2_11_4, n3_11_4);
nor gn5_11_4(n5_11_4, A11B5, n4_11_4);
nor gn6_11_4(n6_11_4, A11B5, n5_11_4);
nor gn7_11_4(n7_11_4, n4_11_4, n5_11_4);
nor gn8_11_4(S11_4, n6_11_4, n7_11_4);
nor gn9_11_4(C11_4, n1_11_4, n5_11_4);

/* FA MFA12_4(S12_4,C12_4,S13_3,C12_3,A12B5); */
nor gn1_12_4(n1_12_4, S13_3, C12_3);
nor gn2_12_4(n2_12_4, n1_12_4, C12_3);
nor gn3_12_4(n3_12_4, S13_3, n1_12_4);
nor gn4_12_4(n4_12_4, n2_12_4, n3_12_4);
nor gn5_12_4(n5_12_4, A12B5, n4_12_4);
nor gn6_12_4(n6_12_4, A12B5, n5_12_4);
nor gn7_12_4(n7_12_4, n4_12_4, n5_12_4);
nor gn8_12_4(S12_4, n6_12_4, n7_12_4);
nor gn9_12_4(C12_4, n1_12_4, n5_12_4);

/* FA MFA13_4(S13_4,C13_4,S14_3,C13_3,A13B5); */
nor gn1_13_4(n1_13_4, S14_3, C13_3);
nor gn2_13_4(n2_13_4, n1_13_4, C13_3);
nor gn3_13_4(n3_13_4, S14_3, n1_13_4);
nor gn4_13_4(n4_13_4, n2_13_4, n3_13_4);
nor gn5_13_4(n5_13_4, A13B5, n4_13_4);
nor gn6_13_4(n6_13_4, A13B5, n5_13_4);
nor gn7_13_4(n7_13_4, n4_13_4, n5_13_4);
nor gn8_13_4(S13_4, n6_13_4, n7_13_4);
nor gn9_13_4(C13_4, n1_13_4, n5_13_4);

/* FA MFA14_4(S14_4,C14_4,A15B4,C14_3,A14B5); */
nor gn1_14_4(n1_14_4, A15B4, C14_3);
nor gn2_14_4(n2_14_4, n1_14_4, C14_3);
nor gn3_14_4(n3_14_4, A15B4, n1_14_4);
nor gn4_14_4(n4_14_4, n2_14_4, n3_14_4);
nor gn5_14_4(n5_14_4, A14B5, n4_14_4);
nor gn6_14_4(n6_14_4, A14B5, n5_14_4);
nor gn7_14_4(n7_14_4, n4_14_4, n5_14_4);
nor gn8_14_4(S14_4, n6_14_4, n7_14_4);
nor gn9_14_4(C14_4, n1_14_4, n5_14_4);

/* FA MFA0_5(S0_5,C0_5,S1_4,C0_4,A0B6); */
nor gn1_0_5(n1_0_5, S1_4, C0_4);
nor gn2_0_5(n2_0_5, n1_0_5, C0_4);
nor gn3_0_5(n3_0_5, S1_4, n1_0_5);
nor gn4_0_5(n4_0_5, n2_0_5, n3_0_5);
nor gn5_0_5(n5_0_5, A0B6, n4_0_5);
nor gn6_0_5(n6_0_5, A0B6, n5_0_5);
nor gn7_0_5(n7_0_5, n4_0_5, n5_0_5);
nor gn8_0_5(S0_5, n6_0_5, n7_0_5);
nor gn9_0_5(C0_5, n1_0_5, n5_0_5);

/* FA MFA1_5(S1_5,C1_5,S2_4,C1_4,A1B6); */
nor gn1_1_5(n1_1_5, S2_4, C1_4);
nor gn2_1_5(n2_1_5, n1_1_5, C1_4);
nor gn3_1_5(n3_1_5, S2_4, n1_1_5);
nor gn4_1_5(n4_1_5, n2_1_5, n3_1_5);
nor gn5_1_5(n5_1_5, A1B6, n4_1_5);
nor gn6_1_5(n6_1_5, A1B6, n5_1_5);
nor gn7_1_5(n7_1_5, n4_1_5, n5_1_5);
nor gn8_1_5(S1_5, n6_1_5, n7_1_5);
nor gn9_1_5(C1_5, n1_1_5, n5_1_5);

/* FA MFA2_5(S2_5,C2_5,S3_4,C2_4,A2B6); */
nor gn1_2_5(n1_2_5, S3_4, C2_4);
nor gn2_2_5(n2_2_5, n1_2_5, C2_4);
nor gn3_2_5(n3_2_5, S3_4, n1_2_5);
nor gn4_2_5(n4_2_5, n2_2_5, n3_2_5);
nor gn5_2_5(n5_2_5, A2B6, n4_2_5);
nor gn6_2_5(n6_2_5, A2B6, n5_2_5);
nor gn7_2_5(n7_2_5, n4_2_5, n5_2_5);
nor gn8_2_5(S2_5, n6_2_5, n7_2_5);
nor gn9_2_5(C2_5, n1_2_5, n5_2_5);

/* FA MFA3_5(S3_5,C3_5,S4_4,C3_4,A3B6); */
nor gn1_3_5(n1_3_5, S4_4, C3_4);
nor gn2_3_5(n2_3_5, n1_3_5, C3_4);
nor gn3_3_5(n3_3_5, S4_4, n1_3_5);
nor gn4_3_5(n4_3_5, n2_3_5, n3_3_5);
nor gn5_3_5(n5_3_5, A3B6, n4_3_5);
nor gn6_3_5(n6_3_5, A3B6, n5_3_5);
nor gn7_3_5(n7_3_5, n4_3_5, n5_3_5);
nor gn8_3_5(S3_5, n6_3_5, n7_3_5);
nor gn9_3_5(C3_5, n1_3_5, n5_3_5);

/* FA MFA4_5(S4_5,C4_5,S5_4,C4_4,A4B6); */
nor gn1_4_5(n1_4_5, S5_4, C4_4);
nor gn2_4_5(n2_4_5, n1_4_5, C4_4);
nor gn3_4_5(n3_4_5, S5_4, n1_4_5);
nor gn4_4_5(n4_4_5, n2_4_5, n3_4_5);
nor gn5_4_5(n5_4_5, A4B6, n4_4_5);
nor gn6_4_5(n6_4_5, A4B6, n5_4_5);
nor gn7_4_5(n7_4_5, n4_4_5, n5_4_5);
nor gn8_4_5(S4_5, n6_4_5, n7_4_5);
nor gn9_4_5(C4_5, n1_4_5, n5_4_5);

/* FA MFA5_5(S5_5,C5_5,S6_4,C5_4,A5B6); */
nor gn1_5_5(n1_5_5, S6_4, C5_4);
nor gn2_5_5(n2_5_5, n1_5_5, C5_4);
nor gn3_5_5(n3_5_5, S6_4, n1_5_5);
nor gn4_5_5(n4_5_5, n2_5_5, n3_5_5);
nor gn5_5_5(n5_5_5, A5B6, n4_5_5);
nor gn6_5_5(n6_5_5, A5B6, n5_5_5);
nor gn7_5_5(n7_5_5, n4_5_5, n5_5_5);
nor gn8_5_5(S5_5, n6_5_5, n7_5_5);
nor gn9_5_5(C5_5, n1_5_5, n5_5_5);

/* FA MFA6_5(S6_5,C6_5,S7_4,C6_4,A6B6); */
nor gn1_6_5(n1_6_5, S7_4, C6_4);
nor gn2_6_5(n2_6_5, n1_6_5, C6_4);
nor gn3_6_5(n3_6_5, S7_4, n1_6_5);
nor gn4_6_5(n4_6_5, n2_6_5, n3_6_5);
nor gn5_6_5(n5_6_5, A6B6, n4_6_5);
nor gn6_6_5(n6_6_5, A6B6, n5_6_5);
nor gn7_6_5(n7_6_5, n4_6_5, n5_6_5);
nor gn8_6_5(S6_5, n6_6_5, n7_6_5);
nor gn9_6_5(C6_5, n1_6_5, n5_6_5);

/* FA MFA7_5(S7_5,C7_5,S8_4,C7_4,A7B6); */
nor gn1_7_5(n1_7_5, S8_4, C7_4);
nor gn2_7_5(n2_7_5, n1_7_5, C7_4);
nor gn3_7_5(n3_7_5, S8_4, n1_7_5);
nor gn4_7_5(n4_7_5, n2_7_5, n3_7_5);
nor gn5_7_5(n5_7_5, A7B6, n4_7_5);
nor gn6_7_5(n6_7_5, A7B6, n5_7_5);
nor gn7_7_5(n7_7_5, n4_7_5, n5_7_5);
nor gn8_7_5(S7_5, n6_7_5, n7_7_5);
nor gn9_7_5(C7_5, n1_7_5, n5_7_5);

/* FA MFA8_5(S8_5,C8_5,S9_4,C8_4,A8B6); */
nor gn1_8_5(n1_8_5, S9_4, C8_4);
nor gn2_8_5(n2_8_5, n1_8_5, C8_4);
nor gn3_8_5(n3_8_5, S9_4, n1_8_5);
nor gn4_8_5(n4_8_5, n2_8_5, n3_8_5);
nor gn5_8_5(n5_8_5, A8B6, n4_8_5);
nor gn6_8_5(n6_8_5, A8B6, n5_8_5);
nor gn7_8_5(n7_8_5, n4_8_5, n5_8_5);
nor gn8_8_5(S8_5, n6_8_5, n7_8_5);
nor gn9_8_5(C8_5, n1_8_5, n5_8_5);

/* FA MFA9_5(S9_5,C9_5,S10_4,C9_4,A9B6); */
nor gn1_9_5(n1_9_5, S10_4, C9_4);
nor gn2_9_5(n2_9_5, n1_9_5, C9_4);
nor gn3_9_5(n3_9_5, S10_4, n1_9_5);
nor gn4_9_5(n4_9_5, n2_9_5, n3_9_5);
nor gn5_9_5(n5_9_5, A9B6, n4_9_5);
nor gn6_9_5(n6_9_5, A9B6, n5_9_5);
nor gn7_9_5(n7_9_5, n4_9_5, n5_9_5);
nor gn8_9_5(S9_5, n6_9_5, n7_9_5);
nor gn9_9_5(C9_5, n1_9_5, n5_9_5);

/* FA MFA10_5(S10_5,C10_5,S11_4,C10_4,A10B6); */
nor gn1_10_5(n1_10_5, S11_4, C10_4);
nor gn2_10_5(n2_10_5, n1_10_5, C10_4);
nor gn3_10_5(n3_10_5, S11_4, n1_10_5);
nor gn4_10_5(n4_10_5, n2_10_5, n3_10_5);
nor gn5_10_5(n5_10_5, A10B6, n4_10_5);
nor gn6_10_5(n6_10_5, A10B6, n5_10_5);
nor gn7_10_5(n7_10_5, n4_10_5, n5_10_5);
nor gn8_10_5(S10_5, n6_10_5, n7_10_5);
nor gn9_10_5(C10_5, n1_10_5, n5_10_5);

/* FA MFA11_5(S11_5,C11_5,S12_4,C11_4,A11B6); */
nor gn1_11_5(n1_11_5, S12_4, C11_4);
nor gn2_11_5(n2_11_5, n1_11_5, C11_4);
nor gn3_11_5(n3_11_5, S12_4, n1_11_5);
nor gn4_11_5(n4_11_5, n2_11_5, n3_11_5);
nor gn5_11_5(n5_11_5, A11B6, n4_11_5);
nor gn6_11_5(n6_11_5, A11B6, n5_11_5);
nor gn7_11_5(n7_11_5, n4_11_5, n5_11_5);
nor gn8_11_5(S11_5, n6_11_5, n7_11_5);
nor gn9_11_5(C11_5, n1_11_5, n5_11_5);

/* FA MFA12_5(S12_5,C12_5,S13_4,C12_4,A12B6); */
nor gn1_12_5(n1_12_5, S13_4, C12_4);
nor gn2_12_5(n2_12_5, n1_12_5, C12_4);
nor gn3_12_5(n3_12_5, S13_4, n1_12_5);
nor gn4_12_5(n4_12_5, n2_12_5, n3_12_5);
nor gn5_12_5(n5_12_5, A12B6, n4_12_5);
nor gn6_12_5(n6_12_5, A12B6, n5_12_5);
nor gn7_12_5(n7_12_5, n4_12_5, n5_12_5);
nor gn8_12_5(S12_5, n6_12_5, n7_12_5);
nor gn9_12_5(C12_5, n1_12_5, n5_12_5);

/* FA MFA13_5(S13_5,C13_5,S14_4,C13_4,A13B6); */
nor gn1_13_5(n1_13_5, S14_4, C13_4);
nor gn2_13_5(n2_13_5, n1_13_5, C13_4);
nor gn3_13_5(n3_13_5, S14_4, n1_13_5);
nor gn4_13_5(n4_13_5, n2_13_5, n3_13_5);
nor gn5_13_5(n5_13_5, A13B6, n4_13_5);
nor gn6_13_5(n6_13_5, A13B6, n5_13_5);
nor gn7_13_5(n7_13_5, n4_13_5, n5_13_5);
nor gn8_13_5(S13_5, n6_13_5, n7_13_5);
nor gn9_13_5(C13_5, n1_13_5, n5_13_5);

/* FA MFA14_5(S14_5,C14_5,A15B5,C14_4,A14B6); */
nor gn1_14_5(n1_14_5, A15B5, C14_4);
nor gn2_14_5(n2_14_5, n1_14_5, C14_4);
nor gn3_14_5(n3_14_5, A15B5, n1_14_5);
nor gn4_14_5(n4_14_5, n2_14_5, n3_14_5);
nor gn5_14_5(n5_14_5, A14B6, n4_14_5);
nor gn6_14_5(n6_14_5, A14B6, n5_14_5);
nor gn7_14_5(n7_14_5, n4_14_5, n5_14_5);
nor gn8_14_5(S14_5, n6_14_5, n7_14_5);
nor gn9_14_5(C14_5, n1_14_5, n5_14_5);

/* FA MFA0_6(S0_6,C0_6,S1_5,C0_5,A0B7); */
nor gn1_0_6(n1_0_6, S1_5, C0_5);
nor gn2_0_6(n2_0_6, n1_0_6, C0_5);
nor gn3_0_6(n3_0_6, S1_5, n1_0_6);
nor gn4_0_6(n4_0_6, n2_0_6, n3_0_6);
nor gn5_0_6(n5_0_6, A0B7, n4_0_6);
nor gn6_0_6(n6_0_6, A0B7, n5_0_6);
nor gn7_0_6(n7_0_6, n4_0_6, n5_0_6);
nor gn8_0_6(S0_6, n6_0_6, n7_0_6);
nor gn9_0_6(C0_6, n1_0_6, n5_0_6);

/* FA MFA1_6(S1_6,C1_6,S2_5,C1_5,A1B7); */
nor gn1_1_6(n1_1_6, S2_5, C1_5);
nor gn2_1_6(n2_1_6, n1_1_6, C1_5);
nor gn3_1_6(n3_1_6, S2_5, n1_1_6);
nor gn4_1_6(n4_1_6, n2_1_6, n3_1_6);
nor gn5_1_6(n5_1_6, A1B7, n4_1_6);
nor gn6_1_6(n6_1_6, A1B7, n5_1_6);
nor gn7_1_6(n7_1_6, n4_1_6, n5_1_6);
nor gn8_1_6(S1_6, n6_1_6, n7_1_6);
nor gn9_1_6(C1_6, n1_1_6, n5_1_6);

/* FA MFA2_6(S2_6,C2_6,S3_5,C2_5,A2B7); */
nor gn1_2_6(n1_2_6, S3_5, C2_5);
nor gn2_2_6(n2_2_6, n1_2_6, C2_5);
nor gn3_2_6(n3_2_6, S3_5, n1_2_6);
nor gn4_2_6(n4_2_6, n2_2_6, n3_2_6);
nor gn5_2_6(n5_2_6, A2B7, n4_2_6);
nor gn6_2_6(n6_2_6, A2B7, n5_2_6);
nor gn7_2_6(n7_2_6, n4_2_6, n5_2_6);
nor gn8_2_6(S2_6, n6_2_6, n7_2_6);
nor gn9_2_6(C2_6, n1_2_6, n5_2_6);

/* FA MFA3_6(S3_6,C3_6,S4_5,C3_5,A3B7); */
nor gn1_3_6(n1_3_6, S4_5, C3_5);
nor gn2_3_6(n2_3_6, n1_3_6, C3_5);
nor gn3_3_6(n3_3_6, S4_5, n1_3_6);
nor gn4_3_6(n4_3_6, n2_3_6, n3_3_6);
nor gn5_3_6(n5_3_6, A3B7, n4_3_6);
nor gn6_3_6(n6_3_6, A3B7, n5_3_6);
nor gn7_3_6(n7_3_6, n4_3_6, n5_3_6);
nor gn8_3_6(S3_6, n6_3_6, n7_3_6);
nor gn9_3_6(C3_6, n1_3_6, n5_3_6);

/* FA MFA4_6(S4_6,C4_6,S5_5,C4_5,A4B7); */
nor gn1_4_6(n1_4_6, S5_5, C4_5);
nor gn2_4_6(n2_4_6, n1_4_6, C4_5);
nor gn3_4_6(n3_4_6, S5_5, n1_4_6);
nor gn4_4_6(n4_4_6, n2_4_6, n3_4_6);
nor gn5_4_6(n5_4_6, A4B7, n4_4_6);
nor gn6_4_6(n6_4_6, A4B7, n5_4_6);
nor gn7_4_6(n7_4_6, n4_4_6, n5_4_6);
nor gn8_4_6(S4_6, n6_4_6, n7_4_6);
nor gn9_4_6(C4_6, n1_4_6, n5_4_6);

/* FA MFA5_6(S5_6,C5_6,S6_5,C5_5,A5B7); */
nor gn1_5_6(n1_5_6, S6_5, C5_5);
nor gn2_5_6(n2_5_6, n1_5_6, C5_5);
nor gn3_5_6(n3_5_6, S6_5, n1_5_6);
nor gn4_5_6(n4_5_6, n2_5_6, n3_5_6);
nor gn5_5_6(n5_5_6, A5B7, n4_5_6);
nor gn6_5_6(n6_5_6, A5B7, n5_5_6);
nor gn7_5_6(n7_5_6, n4_5_6, n5_5_6);
nor gn8_5_6(S5_6, n6_5_6, n7_5_6);
nor gn9_5_6(C5_6, n1_5_6, n5_5_6);

/* FA MFA6_6(S6_6,C6_6,S7_5,C6_5,A6B7); */
nor gn1_6_6(n1_6_6, S7_5, C6_5);
nor gn2_6_6(n2_6_6, n1_6_6, C6_5);
nor gn3_6_6(n3_6_6, S7_5, n1_6_6);
nor gn4_6_6(n4_6_6, n2_6_6, n3_6_6);
nor gn5_6_6(n5_6_6, A6B7, n4_6_6);
nor gn6_6_6(n6_6_6, A6B7, n5_6_6);
nor gn7_6_6(n7_6_6, n4_6_6, n5_6_6);
nor gn8_6_6(S6_6, n6_6_6, n7_6_6);
nor gn9_6_6(C6_6, n1_6_6, n5_6_6);

/* FA MFA7_6(S7_6,C7_6,S8_5,C7_5,A7B7); */
nor gn1_7_6(n1_7_6, S8_5, C7_5);
nor gn2_7_6(n2_7_6, n1_7_6, C7_5);
nor gn3_7_6(n3_7_6, S8_5, n1_7_6);
nor gn4_7_6(n4_7_6, n2_7_6, n3_7_6);
nor gn5_7_6(n5_7_6, A7B7, n4_7_6);
nor gn6_7_6(n6_7_6, A7B7, n5_7_6);
nor gn7_7_6(n7_7_6, n4_7_6, n5_7_6);
nor gn8_7_6(S7_6, n6_7_6, n7_7_6);
nor gn9_7_6(C7_6, n1_7_6, n5_7_6);

/* FA MFA8_6(S8_6,C8_6,S9_5,C8_5,A8B7); */
nor gn1_8_6(n1_8_6, S9_5, C8_5);
nor gn2_8_6(n2_8_6, n1_8_6, C8_5);
nor gn3_8_6(n3_8_6, S9_5, n1_8_6);
nor gn4_8_6(n4_8_6, n2_8_6, n3_8_6);
nor gn5_8_6(n5_8_6, A8B7, n4_8_6);
nor gn6_8_6(n6_8_6, A8B7, n5_8_6);
nor gn7_8_6(n7_8_6, n4_8_6, n5_8_6);
nor gn8_8_6(S8_6, n6_8_6, n7_8_6);
nor gn9_8_6(C8_6, n1_8_6, n5_8_6);

/* FA MFA9_6(S9_6,C9_6,S10_5,C9_5,A9B7); */
nor gn1_9_6(n1_9_6, S10_5, C9_5);
nor gn2_9_6(n2_9_6, n1_9_6, C9_5);
nor gn3_9_6(n3_9_6, S10_5, n1_9_6);
nor gn4_9_6(n4_9_6, n2_9_6, n3_9_6);
nor gn5_9_6(n5_9_6, A9B7, n4_9_6);
nor gn6_9_6(n6_9_6, A9B7, n5_9_6);
nor gn7_9_6(n7_9_6, n4_9_6, n5_9_6);
nor gn8_9_6(S9_6, n6_9_6, n7_9_6);
nor gn9_9_6(C9_6, n1_9_6, n5_9_6);

/* FA MFA10_6(S10_6,C10_6,S11_5,C10_5,A10B7); */
nor gn1_10_6(n1_10_6, S11_5, C10_5);
nor gn2_10_6(n2_10_6, n1_10_6, C10_5);
nor gn3_10_6(n3_10_6, S11_5, n1_10_6);
nor gn4_10_6(n4_10_6, n2_10_6, n3_10_6);
nor gn5_10_6(n5_10_6, A10B7, n4_10_6);
nor gn6_10_6(n6_10_6, A10B7, n5_10_6);
nor gn7_10_6(n7_10_6, n4_10_6, n5_10_6);
nor gn8_10_6(S10_6, n6_10_6, n7_10_6);
nor gn9_10_6(C10_6, n1_10_6, n5_10_6);

/* FA MFA11_6(S11_6,C11_6,S12_5,C11_5,A11B7); */
nor gn1_11_6(n1_11_6, S12_5, C11_5);
nor gn2_11_6(n2_11_6, n1_11_6, C11_5);
nor gn3_11_6(n3_11_6, S12_5, n1_11_6);
nor gn4_11_6(n4_11_6, n2_11_6, n3_11_6);
nor gn5_11_6(n5_11_6, A11B7, n4_11_6);
nor gn6_11_6(n6_11_6, A11B7, n5_11_6);
nor gn7_11_6(n7_11_6, n4_11_6, n5_11_6);
nor gn8_11_6(S11_6, n6_11_6, n7_11_6);
nor gn9_11_6(C11_6, n1_11_6, n5_11_6);

/* FA MFA12_6(S12_6,C12_6,S13_5,C12_5,A12B7); */
nor gn1_12_6(n1_12_6, S13_5, C12_5);
nor gn2_12_6(n2_12_6, n1_12_6, C12_5);
nor gn3_12_6(n3_12_6, S13_5, n1_12_6);
nor gn4_12_6(n4_12_6, n2_12_6, n3_12_6);
nor gn5_12_6(n5_12_6, A12B7, n4_12_6);
nor gn6_12_6(n6_12_6, A12B7, n5_12_6);
nor gn7_12_6(n7_12_6, n4_12_6, n5_12_6);
nor gn8_12_6(S12_6, n6_12_6, n7_12_6);
nor gn9_12_6(C12_6, n1_12_6, n5_12_6);

/* FA MFA13_6(S13_6,C13_6,S14_5,C13_5,A13B7); */
nor gn1_13_6(n1_13_6, S14_5, C13_5);
nor gn2_13_6(n2_13_6, n1_13_6, C13_5);
nor gn3_13_6(n3_13_6, S14_5, n1_13_6);
nor gn4_13_6(n4_13_6, n2_13_6, n3_13_6);
nor gn5_13_6(n5_13_6, A13B7, n4_13_6);
nor gn6_13_6(n6_13_6, A13B7, n5_13_6);
nor gn7_13_6(n7_13_6, n4_13_6, n5_13_6);
nor gn8_13_6(S13_6, n6_13_6, n7_13_6);
nor gn9_13_6(C13_6, n1_13_6, n5_13_6);

/* FA MFA14_6(S14_6,C14_6,A15B6,C14_5,A14B7); */
nor gn1_14_6(n1_14_6, A15B6, C14_5);
nor gn2_14_6(n2_14_6, n1_14_6, C14_5);
nor gn3_14_6(n3_14_6, A15B6, n1_14_6);
nor gn4_14_6(n4_14_6, n2_14_6, n3_14_6);
nor gn5_14_6(n5_14_6, A14B7, n4_14_6);
nor gn6_14_6(n6_14_6, A14B7, n5_14_6);
nor gn7_14_6(n7_14_6, n4_14_6, n5_14_6);
nor gn8_14_6(S14_6, n6_14_6, n7_14_6);
nor gn9_14_6(C14_6, n1_14_6, n5_14_6);

/* FA MFA0_7(S0_7,C0_7,S1_6,C0_6,A0B8); */
nor gn1_0_7(n1_0_7, S1_6, C0_6);
nor gn2_0_7(n2_0_7, n1_0_7, C0_6);
nor gn3_0_7(n3_0_7, S1_6, n1_0_7);
nor gn4_0_7(n4_0_7, n2_0_7, n3_0_7);
nor gn5_0_7(n5_0_7, A0B8, n4_0_7);
nor gn6_0_7(n6_0_7, A0B8, n5_0_7);
nor gn7_0_7(n7_0_7, n4_0_7, n5_0_7);
nor gn8_0_7(S0_7, n6_0_7, n7_0_7);
nor gn9_0_7(C0_7, n1_0_7, n5_0_7);

/* FA MFA1_7(S1_7,C1_7,S2_6,C1_6,A1B8); */
nor gn1_1_7(n1_1_7, S2_6, C1_6);
nor gn2_1_7(n2_1_7, n1_1_7, C1_6);
nor gn3_1_7(n3_1_7, S2_6, n1_1_7);
nor gn4_1_7(n4_1_7, n2_1_7, n3_1_7);
nor gn5_1_7(n5_1_7, A1B8, n4_1_7);
nor gn6_1_7(n6_1_7, A1B8, n5_1_7);
nor gn7_1_7(n7_1_7, n4_1_7, n5_1_7);
nor gn8_1_7(S1_7, n6_1_7, n7_1_7);
nor gn9_1_7(C1_7, n1_1_7, n5_1_7);

/* FA MFA2_7(S2_7,C2_7,S3_6,C2_6,A2B8); */
nor gn1_2_7(n1_2_7, S3_6, C2_6);
nor gn2_2_7(n2_2_7, n1_2_7, C2_6);
nor gn3_2_7(n3_2_7, S3_6, n1_2_7);
nor gn4_2_7(n4_2_7, n2_2_7, n3_2_7);
nor gn5_2_7(n5_2_7, A2B8, n4_2_7);
nor gn6_2_7(n6_2_7, A2B8, n5_2_7);
nor gn7_2_7(n7_2_7, n4_2_7, n5_2_7);
nor gn8_2_7(S2_7, n6_2_7, n7_2_7);
nor gn9_2_7(C2_7, n1_2_7, n5_2_7);

/* FA MFA3_7(S3_7,C3_7,S4_6,C3_6,A3B8); */
nor gn1_3_7(n1_3_7, S4_6, C3_6);
nor gn2_3_7(n2_3_7, n1_3_7, C3_6);
nor gn3_3_7(n3_3_7, S4_6, n1_3_7);
nor gn4_3_7(n4_3_7, n2_3_7, n3_3_7);
nor gn5_3_7(n5_3_7, A3B8, n4_3_7);
nor gn6_3_7(n6_3_7, A3B8, n5_3_7);
nor gn7_3_7(n7_3_7, n4_3_7, n5_3_7);
nor gn8_3_7(S3_7, n6_3_7, n7_3_7);
nor gn9_3_7(C3_7, n1_3_7, n5_3_7);

/* FA MFA4_7(S4_7,C4_7,S5_6,C4_6,A4B8); */
nor gn1_4_7(n1_4_7, S5_6, C4_6);
nor gn2_4_7(n2_4_7, n1_4_7, C4_6);
nor gn3_4_7(n3_4_7, S5_6, n1_4_7);
nor gn4_4_7(n4_4_7, n2_4_7, n3_4_7);
nor gn5_4_7(n5_4_7, A4B8, n4_4_7);
nor gn6_4_7(n6_4_7, A4B8, n5_4_7);
nor gn7_4_7(n7_4_7, n4_4_7, n5_4_7);
nor gn8_4_7(S4_7, n6_4_7, n7_4_7);
nor gn9_4_7(C4_7, n1_4_7, n5_4_7);

/* FA MFA5_7(S5_7,C5_7,S6_6,C5_6,A5B8); */
nor gn1_5_7(n1_5_7, S6_6, C5_6);
nor gn2_5_7(n2_5_7, n1_5_7, C5_6);
nor gn3_5_7(n3_5_7, S6_6, n1_5_7);
nor gn4_5_7(n4_5_7, n2_5_7, n3_5_7);
nor gn5_5_7(n5_5_7, A5B8, n4_5_7);
nor gn6_5_7(n6_5_7, A5B8, n5_5_7);
nor gn7_5_7(n7_5_7, n4_5_7, n5_5_7);
nor gn8_5_7(S5_7, n6_5_7, n7_5_7);
nor gn9_5_7(C5_7, n1_5_7, n5_5_7);

/* FA MFA6_7(S6_7,C6_7,S7_6,C6_6,A6B8); */
nor gn1_6_7(n1_6_7, S7_6, C6_6);
nor gn2_6_7(n2_6_7, n1_6_7, C6_6);
nor gn3_6_7(n3_6_7, S7_6, n1_6_7);
nor gn4_6_7(n4_6_7, n2_6_7, n3_6_7);
nor gn5_6_7(n5_6_7, A6B8, n4_6_7);
nor gn6_6_7(n6_6_7, A6B8, n5_6_7);
nor gn7_6_7(n7_6_7, n4_6_7, n5_6_7);
nor gn8_6_7(S6_7, n6_6_7, n7_6_7);
nor gn9_6_7(C6_7, n1_6_7, n5_6_7);

/* FA MFA7_7(S7_7,C7_7,S8_6,C7_6,A7B8); */
nor gn1_7_7(n1_7_7, S8_6, C7_6);
nor gn2_7_7(n2_7_7, n1_7_7, C7_6);
nor gn3_7_7(n3_7_7, S8_6, n1_7_7);
nor gn4_7_7(n4_7_7, n2_7_7, n3_7_7);
nor gn5_7_7(n5_7_7, A7B8, n4_7_7);
nor gn6_7_7(n6_7_7, A7B8, n5_7_7);
nor gn7_7_7(n7_7_7, n4_7_7, n5_7_7);
nor gn8_7_7(S7_7, n6_7_7, n7_7_7);
nor gn9_7_7(C7_7, n1_7_7, n5_7_7);

/* FA MFA8_7(S8_7,C8_7,S9_6,C8_6,A8B8); */
nor gn1_8_7(n1_8_7, S9_6, C8_6);
nor gn2_8_7(n2_8_7, n1_8_7, C8_6);
nor gn3_8_7(n3_8_7, S9_6, n1_8_7);
nor gn4_8_7(n4_8_7, n2_8_7, n3_8_7);
nor gn5_8_7(n5_8_7, A8B8, n4_8_7);
nor gn6_8_7(n6_8_7, A8B8, n5_8_7);
nor gn7_8_7(n7_8_7, n4_8_7, n5_8_7);
nor gn8_8_7(S8_7, n6_8_7, n7_8_7);
nor gn9_8_7(C8_7, n1_8_7, n5_8_7);

/* FA MFA9_7(S9_7,C9_7,S10_6,C9_6,A9B8); */
nor gn1_9_7(n1_9_7, S10_6, C9_6);
nor gn2_9_7(n2_9_7, n1_9_7, C9_6);
nor gn3_9_7(n3_9_7, S10_6, n1_9_7);
nor gn4_9_7(n4_9_7, n2_9_7, n3_9_7);
nor gn5_9_7(n5_9_7, A9B8, n4_9_7);
nor gn6_9_7(n6_9_7, A9B8, n5_9_7);
nor gn7_9_7(n7_9_7, n4_9_7, n5_9_7);
nor gn8_9_7(S9_7, n6_9_7, n7_9_7);
nor gn9_9_7(C9_7, n1_9_7, n5_9_7);

/* FA MFA10_7(S10_7,C10_7,S11_6,C10_6,A10B8); */
nor gn1_10_7(n1_10_7, S11_6, C10_6);
nor gn2_10_7(n2_10_7, n1_10_7, C10_6);
nor gn3_10_7(n3_10_7, S11_6, n1_10_7);
nor gn4_10_7(n4_10_7, n2_10_7, n3_10_7);
nor gn5_10_7(n5_10_7, A10B8, n4_10_7);
nor gn6_10_7(n6_10_7, A10B8, n5_10_7);
nor gn7_10_7(n7_10_7, n4_10_7, n5_10_7);
nor gn8_10_7(S10_7, n6_10_7, n7_10_7);
nor gn9_10_7(C10_7, n1_10_7, n5_10_7);

/* FA MFA11_7(S11_7,C11_7,S12_6,C11_6,A11B8); */
nor gn1_11_7(n1_11_7, S12_6, C11_6);
nor gn2_11_7(n2_11_7, n1_11_7, C11_6);
nor gn3_11_7(n3_11_7, S12_6, n1_11_7);
nor gn4_11_7(n4_11_7, n2_11_7, n3_11_7);
nor gn5_11_7(n5_11_7, A11B8, n4_11_7);
nor gn6_11_7(n6_11_7, A11B8, n5_11_7);
nor gn7_11_7(n7_11_7, n4_11_7, n5_11_7);
nor gn8_11_7(S11_7, n6_11_7, n7_11_7);
nor gn9_11_7(C11_7, n1_11_7, n5_11_7);

/* FA MFA12_7(S12_7,C12_7,S13_6,C12_6,A12B8); */
nor gn1_12_7(n1_12_7, S13_6, C12_6);
nor gn2_12_7(n2_12_7, n1_12_7, C12_6);
nor gn3_12_7(n3_12_7, S13_6, n1_12_7);
nor gn4_12_7(n4_12_7, n2_12_7, n3_12_7);
nor gn5_12_7(n5_12_7, A12B8, n4_12_7);
nor gn6_12_7(n6_12_7, A12B8, n5_12_7);
nor gn7_12_7(n7_12_7, n4_12_7, n5_12_7);
nor gn8_12_7(S12_7, n6_12_7, n7_12_7);
nor gn9_12_7(C12_7, n1_12_7, n5_12_7);

/* FA MFA13_7(S13_7,C13_7,S14_6,C13_6,A13B8); */
nor gn1_13_7(n1_13_7, S14_6, C13_6);
nor gn2_13_7(n2_13_7, n1_13_7, C13_6);
nor gn3_13_7(n3_13_7, S14_6, n1_13_7);
nor gn4_13_7(n4_13_7, n2_13_7, n3_13_7);
nor gn5_13_7(n5_13_7, A13B8, n4_13_7);
nor gn6_13_7(n6_13_7, A13B8, n5_13_7);
nor gn7_13_7(n7_13_7, n4_13_7, n5_13_7);
nor gn8_13_7(S13_7, n6_13_7, n7_13_7);
nor gn9_13_7(C13_7, n1_13_7, n5_13_7);

/* FA MFA14_7(S14_7,C14_7,A15B7,C14_6,A14B8); */
nor gn1_14_7(n1_14_7, A15B7, C14_6);
nor gn2_14_7(n2_14_7, n1_14_7, C14_6);
nor gn3_14_7(n3_14_7, A15B7, n1_14_7);
nor gn4_14_7(n4_14_7, n2_14_7, n3_14_7);
nor gn5_14_7(n5_14_7, A14B8, n4_14_7);
nor gn6_14_7(n6_14_7, A14B8, n5_14_7);
nor gn7_14_7(n7_14_7, n4_14_7, n5_14_7);
nor gn8_14_7(S14_7, n6_14_7, n7_14_7);
nor gn9_14_7(C14_7, n1_14_7, n5_14_7);

/* FA MFA0_8(S0_8,C0_8,S1_7,C0_7,A0B9); */
nor gn1_0_8(n1_0_8, S1_7, C0_7);
nor gn2_0_8(n2_0_8, n1_0_8, C0_7);
nor gn3_0_8(n3_0_8, S1_7, n1_0_8);
nor gn4_0_8(n4_0_8, n2_0_8, n3_0_8);
nor gn5_0_8(n5_0_8, A0B9, n4_0_8);
nor gn6_0_8(n6_0_8, A0B9, n5_0_8);
nor gn7_0_8(n7_0_8, n4_0_8, n5_0_8);
nor gn8_0_8(S0_8, n6_0_8, n7_0_8);
nor gn9_0_8(C0_8, n1_0_8, n5_0_8);

/* FA MFA1_8(S1_8,C1_8,S2_7,C1_7,A1B9); */
nor gn1_1_8(n1_1_8, S2_7, C1_7);
nor gn2_1_8(n2_1_8, n1_1_8, C1_7);
nor gn3_1_8(n3_1_8, S2_7, n1_1_8);
nor gn4_1_8(n4_1_8, n2_1_8, n3_1_8);
nor gn5_1_8(n5_1_8, A1B9, n4_1_8);
nor gn6_1_8(n6_1_8, A1B9, n5_1_8);
nor gn7_1_8(n7_1_8, n4_1_8, n5_1_8);
nor gn8_1_8(S1_8, n6_1_8, n7_1_8);
nor gn9_1_8(C1_8, n1_1_8, n5_1_8);

/* FA MFA2_8(S2_8,C2_8,S3_7,C2_7,A2B9); */
nor gn1_2_8(n1_2_8, S3_7, C2_7);
nor gn2_2_8(n2_2_8, n1_2_8, C2_7);
nor gn3_2_8(n3_2_8, S3_7, n1_2_8);
nor gn4_2_8(n4_2_8, n2_2_8, n3_2_8);
nor gn5_2_8(n5_2_8, A2B9, n4_2_8);
nor gn6_2_8(n6_2_8, A2B9, n5_2_8);
nor gn7_2_8(n7_2_8, n4_2_8, n5_2_8);
nor gn8_2_8(S2_8, n6_2_8, n7_2_8);
nor gn9_2_8(C2_8, n1_2_8, n5_2_8);

/* FA MFA3_8(S3_8,C3_8,S4_7,C3_7,A3B9); */
nor gn1_3_8(n1_3_8, S4_7, C3_7);
nor gn2_3_8(n2_3_8, n1_3_8, C3_7);
nor gn3_3_8(n3_3_8, S4_7, n1_3_8);
nor gn4_3_8(n4_3_8, n2_3_8, n3_3_8);
nor gn5_3_8(n5_3_8, A3B9, n4_3_8);
nor gn6_3_8(n6_3_8, A3B9, n5_3_8);
nor gn7_3_8(n7_3_8, n4_3_8, n5_3_8);
nor gn8_3_8(S3_8, n6_3_8, n7_3_8);
nor gn9_3_8(C3_8, n1_3_8, n5_3_8);

/* FA MFA4_8(S4_8,C4_8,S5_7,C4_7,A4B9); */
nor gn1_4_8(n1_4_8, S5_7, C4_7);
nor gn2_4_8(n2_4_8, n1_4_8, C4_7);
nor gn3_4_8(n3_4_8, S5_7, n1_4_8);
nor gn4_4_8(n4_4_8, n2_4_8, n3_4_8);
nor gn5_4_8(n5_4_8, A4B9, n4_4_8);
nor gn6_4_8(n6_4_8, A4B9, n5_4_8);
nor gn7_4_8(n7_4_8, n4_4_8, n5_4_8);
nor gn8_4_8(S4_8, n6_4_8, n7_4_8);
nor gn9_4_8(C4_8, n1_4_8, n5_4_8);

/* FA MFA5_8(S5_8,C5_8,S6_7,C5_7,A5B9); */
nor gn1_5_8(n1_5_8, S6_7, C5_7);
nor gn2_5_8(n2_5_8, n1_5_8, C5_7);
nor gn3_5_8(n3_5_8, S6_7, n1_5_8);
nor gn4_5_8(n4_5_8, n2_5_8, n3_5_8);
nor gn5_5_8(n5_5_8, A5B9, n4_5_8);
nor gn6_5_8(n6_5_8, A5B9, n5_5_8);
nor gn7_5_8(n7_5_8, n4_5_8, n5_5_8);
nor gn8_5_8(S5_8, n6_5_8, n7_5_8);
nor gn9_5_8(C5_8, n1_5_8, n5_5_8);

/* FA MFA6_8(S6_8,C6_8,S7_7,C6_7,A6B9); */
nor gn1_6_8(n1_6_8, S7_7, C6_7);
nor gn2_6_8(n2_6_8, n1_6_8, C6_7);
nor gn3_6_8(n3_6_8, S7_7, n1_6_8);
nor gn4_6_8(n4_6_8, n2_6_8, n3_6_8);
nor gn5_6_8(n5_6_8, A6B9, n4_6_8);
nor gn6_6_8(n6_6_8, A6B9, n5_6_8);
nor gn7_6_8(n7_6_8, n4_6_8, n5_6_8);
nor gn8_6_8(S6_8, n6_6_8, n7_6_8);
nor gn9_6_8(C6_8, n1_6_8, n5_6_8);

/* FA MFA7_8(S7_8,C7_8,S8_7,C7_7,A7B9); */
nor gn1_7_8(n1_7_8, S8_7, C7_7);
nor gn2_7_8(n2_7_8, n1_7_8, C7_7);
nor gn3_7_8(n3_7_8, S8_7, n1_7_8);
nor gn4_7_8(n4_7_8, n2_7_8, n3_7_8);
nor gn5_7_8(n5_7_8, A7B9, n4_7_8);
nor gn6_7_8(n6_7_8, A7B9, n5_7_8);
nor gn7_7_8(n7_7_8, n4_7_8, n5_7_8);
nor gn8_7_8(S7_8, n6_7_8, n7_7_8);
nor gn9_7_8(C7_8, n1_7_8, n5_7_8);

/* FA MFA8_8(S8_8,C8_8,S9_7,C8_7,A8B9); */
nor gn1_8_8(n1_8_8, S9_7, C8_7);
nor gn2_8_8(n2_8_8, n1_8_8, C8_7);
nor gn3_8_8(n3_8_8, S9_7, n1_8_8);
nor gn4_8_8(n4_8_8, n2_8_8, n3_8_8);
nor gn5_8_8(n5_8_8, A8B9, n4_8_8);
nor gn6_8_8(n6_8_8, A8B9, n5_8_8);
nor gn7_8_8(n7_8_8, n4_8_8, n5_8_8);
nor gn8_8_8(S8_8, n6_8_8, n7_8_8);
nor gn9_8_8(C8_8, n1_8_8, n5_8_8);

/* FA MFA9_8(S9_8,C9_8,S10_7,C9_7,A9B9); */
nor gn1_9_8(n1_9_8, S10_7, C9_7);
nor gn2_9_8(n2_9_8, n1_9_8, C9_7);
nor gn3_9_8(n3_9_8, S10_7, n1_9_8);
nor gn4_9_8(n4_9_8, n2_9_8, n3_9_8);
nor gn5_9_8(n5_9_8, A9B9, n4_9_8);
nor gn6_9_8(n6_9_8, A9B9, n5_9_8);
nor gn7_9_8(n7_9_8, n4_9_8, n5_9_8);
nor gn8_9_8(S9_8, n6_9_8, n7_9_8);
nor gn9_9_8(C9_8, n1_9_8, n5_9_8);

/* FA MFA10_8(S10_8,C10_8,S11_7,C10_7,A10B9); */
nor gn1_10_8(n1_10_8, S11_7, C10_7);
nor gn2_10_8(n2_10_8, n1_10_8, C10_7);
nor gn3_10_8(n3_10_8, S11_7, n1_10_8);
nor gn4_10_8(n4_10_8, n2_10_8, n3_10_8);
nor gn5_10_8(n5_10_8, A10B9, n4_10_8);
nor gn6_10_8(n6_10_8, A10B9, n5_10_8);
nor gn7_10_8(n7_10_8, n4_10_8, n5_10_8);
nor gn8_10_8(S10_8, n6_10_8, n7_10_8);
nor gn9_10_8(C10_8, n1_10_8, n5_10_8);

/* FA MFA11_8(S11_8,C11_8,S12_7,C11_7,A11B9); */
nor gn1_11_8(n1_11_8, S12_7, C11_7);
nor gn2_11_8(n2_11_8, n1_11_8, C11_7);
nor gn3_11_8(n3_11_8, S12_7, n1_11_8);
nor gn4_11_8(n4_11_8, n2_11_8, n3_11_8);
nor gn5_11_8(n5_11_8, A11B9, n4_11_8);
nor gn6_11_8(n6_11_8, A11B9, n5_11_8);
nor gn7_11_8(n7_11_8, n4_11_8, n5_11_8);
nor gn8_11_8(S11_8, n6_11_8, n7_11_8);
nor gn9_11_8(C11_8, n1_11_8, n5_11_8);

/* FA MFA12_8(S12_8,C12_8,S13_7,C12_7,A12B9); */
nor gn1_12_8(n1_12_8, S13_7, C12_7);
nor gn2_12_8(n2_12_8, n1_12_8, C12_7);
nor gn3_12_8(n3_12_8, S13_7, n1_12_8);
nor gn4_12_8(n4_12_8, n2_12_8, n3_12_8);
nor gn5_12_8(n5_12_8, A12B9, n4_12_8);
nor gn6_12_8(n6_12_8, A12B9, n5_12_8);
nor gn7_12_8(n7_12_8, n4_12_8, n5_12_8);
nor gn8_12_8(S12_8, n6_12_8, n7_12_8);
nor gn9_12_8(C12_8, n1_12_8, n5_12_8);

/* FA MFA13_8(S13_8,C13_8,S14_7,C13_7,A13B9); */
nor gn1_13_8(n1_13_8, S14_7, C13_7);
nor gn2_13_8(n2_13_8, n1_13_8, C13_7);
nor gn3_13_8(n3_13_8, S14_7, n1_13_8);
nor gn4_13_8(n4_13_8, n2_13_8, n3_13_8);
nor gn5_13_8(n5_13_8, A13B9, n4_13_8);
nor gn6_13_8(n6_13_8, A13B9, n5_13_8);
nor gn7_13_8(n7_13_8, n4_13_8, n5_13_8);
nor gn8_13_8(S13_8, n6_13_8, n7_13_8);
nor gn9_13_8(C13_8, n1_13_8, n5_13_8);

/* FA MFA14_8(S14_8,C14_8,A15B8,C14_7,A14B9); */
nor gn1_14_8(n1_14_8, A15B8, C14_7);
nor gn2_14_8(n2_14_8, n1_14_8, C14_7);
nor gn3_14_8(n3_14_8, A15B8, n1_14_8);
nor gn4_14_8(n4_14_8, n2_14_8, n3_14_8);
nor gn5_14_8(n5_14_8, A14B9, n4_14_8);
nor gn6_14_8(n6_14_8, A14B9, n5_14_8);
nor gn7_14_8(n7_14_8, n4_14_8, n5_14_8);
nor gn8_14_8(S14_8, n6_14_8, n7_14_8);
nor gn9_14_8(C14_8, n1_14_8, n5_14_8);

/* FA MFA0_9(S0_9,C0_9,S1_8,C0_8,A0B10); */
nor gn1_0_9(n1_0_9, S1_8, C0_8);
nor gn2_0_9(n2_0_9, n1_0_9, C0_8);
nor gn3_0_9(n3_0_9, S1_8, n1_0_9);
nor gn4_0_9(n4_0_9, n2_0_9, n3_0_9);
nor gn5_0_9(n5_0_9, A0B10, n4_0_9);
nor gn6_0_9(n6_0_9, A0B10, n5_0_9);
nor gn7_0_9(n7_0_9, n4_0_9, n5_0_9);
nor gn8_0_9(S0_9, n6_0_9, n7_0_9);
nor gn9_0_9(C0_9, n1_0_9, n5_0_9);

/* FA MFA1_9(S1_9,C1_9,S2_8,C1_8,A1B10); */
nor gn1_1_9(n1_1_9, S2_8, C1_8);
nor gn2_1_9(n2_1_9, n1_1_9, C1_8);
nor gn3_1_9(n3_1_9, S2_8, n1_1_9);
nor gn4_1_9(n4_1_9, n2_1_9, n3_1_9);
nor gn5_1_9(n5_1_9, A1B10, n4_1_9);
nor gn6_1_9(n6_1_9, A1B10, n5_1_9);
nor gn7_1_9(n7_1_9, n4_1_9, n5_1_9);
nor gn8_1_9(S1_9, n6_1_9, n7_1_9);
nor gn9_1_9(C1_9, n1_1_9, n5_1_9);

/* FA MFA2_9(S2_9,C2_9,S3_8,C2_8,A2B10); */
nor gn1_2_9(n1_2_9, S3_8, C2_8);
nor gn2_2_9(n2_2_9, n1_2_9, C2_8);
nor gn3_2_9(n3_2_9, S3_8, n1_2_9);
nor gn4_2_9(n4_2_9, n2_2_9, n3_2_9);
nor gn5_2_9(n5_2_9, A2B10, n4_2_9);
nor gn6_2_9(n6_2_9, A2B10, n5_2_9);
nor gn7_2_9(n7_2_9, n4_2_9, n5_2_9);
nor gn8_2_9(S2_9, n6_2_9, n7_2_9);
nor gn9_2_9(C2_9, n1_2_9, n5_2_9);

/* FA MFA3_9(S3_9,C3_9,S4_8,C3_8,A3B10); */
nor gn1_3_9(n1_3_9, S4_8, C3_8);
nor gn2_3_9(n2_3_9, n1_3_9, C3_8);
nor gn3_3_9(n3_3_9, S4_8, n1_3_9);
nor gn4_3_9(n4_3_9, n2_3_9, n3_3_9);
nor gn5_3_9(n5_3_9, A3B10, n4_3_9);
nor gn6_3_9(n6_3_9, A3B10, n5_3_9);
nor gn7_3_9(n7_3_9, n4_3_9, n5_3_9);
nor gn8_3_9(S3_9, n6_3_9, n7_3_9);
nor gn9_3_9(C3_9, n1_3_9, n5_3_9);

/* FA MFA4_9(S4_9,C4_9,S5_8,C4_8,A4B10); */
nor gn1_4_9(n1_4_9, S5_8, C4_8);
nor gn2_4_9(n2_4_9, n1_4_9, C4_8);
nor gn3_4_9(n3_4_9, S5_8, n1_4_9);
nor gn4_4_9(n4_4_9, n2_4_9, n3_4_9);
nor gn5_4_9(n5_4_9, A4B10, n4_4_9);
nor gn6_4_9(n6_4_9, A4B10, n5_4_9);
nor gn7_4_9(n7_4_9, n4_4_9, n5_4_9);
nor gn8_4_9(S4_9, n6_4_9, n7_4_9);
nor gn9_4_9(C4_9, n1_4_9, n5_4_9);

/* FA MFA5_9(S5_9,C5_9,S6_8,C5_8,A5B10); */
nor gn1_5_9(n1_5_9, S6_8, C5_8);
nor gn2_5_9(n2_5_9, n1_5_9, C5_8);
nor gn3_5_9(n3_5_9, S6_8, n1_5_9);
nor gn4_5_9(n4_5_9, n2_5_9, n3_5_9);
nor gn5_5_9(n5_5_9, A5B10, n4_5_9);
nor gn6_5_9(n6_5_9, A5B10, n5_5_9);
nor gn7_5_9(n7_5_9, n4_5_9, n5_5_9);
nor gn8_5_9(S5_9, n6_5_9, n7_5_9);
nor gn9_5_9(C5_9, n1_5_9, n5_5_9);

/* FA MFA6_9(S6_9,C6_9,S7_8,C6_8,A6B10); */
nor gn1_6_9(n1_6_9, S7_8, C6_8);
nor gn2_6_9(n2_6_9, n1_6_9, C6_8);
nor gn3_6_9(n3_6_9, S7_8, n1_6_9);
nor gn4_6_9(n4_6_9, n2_6_9, n3_6_9);
nor gn5_6_9(n5_6_9, A6B10, n4_6_9);
nor gn6_6_9(n6_6_9, A6B10, n5_6_9);
nor gn7_6_9(n7_6_9, n4_6_9, n5_6_9);
nor gn8_6_9(S6_9, n6_6_9, n7_6_9);
nor gn9_6_9(C6_9, n1_6_9, n5_6_9);

/* FA MFA7_9(S7_9,C7_9,S8_8,C7_8,A7B10); */
nor gn1_7_9(n1_7_9, S8_8, C7_8);
nor gn2_7_9(n2_7_9, n1_7_9, C7_8);
nor gn3_7_9(n3_7_9, S8_8, n1_7_9);
nor gn4_7_9(n4_7_9, n2_7_9, n3_7_9);
nor gn5_7_9(n5_7_9, A7B10, n4_7_9);
nor gn6_7_9(n6_7_9, A7B10, n5_7_9);
nor gn7_7_9(n7_7_9, n4_7_9, n5_7_9);
nor gn8_7_9(S7_9, n6_7_9, n7_7_9);
nor gn9_7_9(C7_9, n1_7_9, n5_7_9);

/* FA MFA8_9(S8_9,C8_9,S9_8,C8_8,A8B10); */
nor gn1_8_9(n1_8_9, S9_8, C8_8);
nor gn2_8_9(n2_8_9, n1_8_9, C8_8);
nor gn3_8_9(n3_8_9, S9_8, n1_8_9);
nor gn4_8_9(n4_8_9, n2_8_9, n3_8_9);
nor gn5_8_9(n5_8_9, A8B10, n4_8_9);
nor gn6_8_9(n6_8_9, A8B10, n5_8_9);
nor gn7_8_9(n7_8_9, n4_8_9, n5_8_9);
nor gn8_8_9(S8_9, n6_8_9, n7_8_9);
nor gn9_8_9(C8_9, n1_8_9, n5_8_9);

/* FA MFA9_9(S9_9,C9_9,S10_8,C9_8,A9B10); */
nor gn1_9_9(n1_9_9, S10_8, C9_8);
nor gn2_9_9(n2_9_9, n1_9_9, C9_8);
nor gn3_9_9(n3_9_9, S10_8, n1_9_9);
nor gn4_9_9(n4_9_9, n2_9_9, n3_9_9);
nor gn5_9_9(n5_9_9, A9B10, n4_9_9);
nor gn6_9_9(n6_9_9, A9B10, n5_9_9);
nor gn7_9_9(n7_9_9, n4_9_9, n5_9_9);
nor gn8_9_9(S9_9, n6_9_9, n7_9_9);
nor gn9_9_9(C9_9, n1_9_9, n5_9_9);

/* FA MFA10_9(S10_9,C10_9,S11_8,C10_8,A10B10); */
nor gn1_10_9(n1_10_9, S11_8, C10_8);
nor gn2_10_9(n2_10_9, n1_10_9, C10_8);
nor gn3_10_9(n3_10_9, S11_8, n1_10_9);
nor gn4_10_9(n4_10_9, n2_10_9, n3_10_9);
nor gn5_10_9(n5_10_9, A10B10, n4_10_9);
nor gn6_10_9(n6_10_9, A10B10, n5_10_9);
nor gn7_10_9(n7_10_9, n4_10_9, n5_10_9);
nor gn8_10_9(S10_9, n6_10_9, n7_10_9);
nor gn9_10_9(C10_9, n1_10_9, n5_10_9);

/* FA MFA11_9(S11_9,C11_9,S12_8,C11_8,A11B10); */
nor gn1_11_9(n1_11_9, S12_8, C11_8);
nor gn2_11_9(n2_11_9, n1_11_9, C11_8);
nor gn3_11_9(n3_11_9, S12_8, n1_11_9);
nor gn4_11_9(n4_11_9, n2_11_9, n3_11_9);
nor gn5_11_9(n5_11_9, A11B10, n4_11_9);
nor gn6_11_9(n6_11_9, A11B10, n5_11_9);
nor gn7_11_9(n7_11_9, n4_11_9, n5_11_9);
nor gn8_11_9(S11_9, n6_11_9, n7_11_9);
nor gn9_11_9(C11_9, n1_11_9, n5_11_9);

/* FA MFA12_9(S12_9,C12_9,S13_8,C12_8,A12B10); */
nor gn1_12_9(n1_12_9, S13_8, C12_8);
nor gn2_12_9(n2_12_9, n1_12_9, C12_8);
nor gn3_12_9(n3_12_9, S13_8, n1_12_9);
nor gn4_12_9(n4_12_9, n2_12_9, n3_12_9);
nor gn5_12_9(n5_12_9, A12B10, n4_12_9);
nor gn6_12_9(n6_12_9, A12B10, n5_12_9);
nor gn7_12_9(n7_12_9, n4_12_9, n5_12_9);
nor gn8_12_9(S12_9, n6_12_9, n7_12_9);
nor gn9_12_9(C12_9, n1_12_9, n5_12_9);

/* FA MFA13_9(S13_9,C13_9,S14_8,C13_8,A13B10); */
nor gn1_13_9(n1_13_9, S14_8, C13_8);
nor gn2_13_9(n2_13_9, n1_13_9, C13_8);
nor gn3_13_9(n3_13_9, S14_8, n1_13_9);
nor gn4_13_9(n4_13_9, n2_13_9, n3_13_9);
nor gn5_13_9(n5_13_9, A13B10, n4_13_9);
nor gn6_13_9(n6_13_9, A13B10, n5_13_9);
nor gn7_13_9(n7_13_9, n4_13_9, n5_13_9);
nor gn8_13_9(S13_9, n6_13_9, n7_13_9);
nor gn9_13_9(C13_9, n1_13_9, n5_13_9);

/* FA MFA14_9(S14_9,C14_9,A15B9,C14_8,A14B10); */
nor gn1_14_9(n1_14_9, A15B9, C14_8);
nor gn2_14_9(n2_14_9, n1_14_9, C14_8);
nor gn3_14_9(n3_14_9, A15B9, n1_14_9);
nor gn4_14_9(n4_14_9, n2_14_9, n3_14_9);
nor gn5_14_9(n5_14_9, A14B10, n4_14_9);
nor gn6_14_9(n6_14_9, A14B10, n5_14_9);
nor gn7_14_9(n7_14_9, n4_14_9, n5_14_9);
nor gn8_14_9(S14_9, n6_14_9, n7_14_9);
nor gn9_14_9(C14_9, n1_14_9, n5_14_9);

/* FA MFA0_10(S0_10,C0_10,S1_9,C0_9,A0B11); */
nor gn1_0_10(n1_0_10, S1_9, C0_9);
nor gn2_0_10(n2_0_10, n1_0_10, C0_9);
nor gn3_0_10(n3_0_10, S1_9, n1_0_10);
nor gn4_0_10(n4_0_10, n2_0_10, n3_0_10);
nor gn5_0_10(n5_0_10, A0B11, n4_0_10);
nor gn6_0_10(n6_0_10, A0B11, n5_0_10);
nor gn7_0_10(n7_0_10, n4_0_10, n5_0_10);
nor gn8_0_10(S0_10, n6_0_10, n7_0_10);
nor gn9_0_10(C0_10, n1_0_10, n5_0_10);

/* FA MFA1_10(S1_10,C1_10,S2_9,C1_9,A1B11); */
nor gn1_1_10(n1_1_10, S2_9, C1_9);
nor gn2_1_10(n2_1_10, n1_1_10, C1_9);
nor gn3_1_10(n3_1_10, S2_9, n1_1_10);
nor gn4_1_10(n4_1_10, n2_1_10, n3_1_10);
nor gn5_1_10(n5_1_10, A1B11, n4_1_10);
nor gn6_1_10(n6_1_10, A1B11, n5_1_10);
nor gn7_1_10(n7_1_10, n4_1_10, n5_1_10);
nor gn8_1_10(S1_10, n6_1_10, n7_1_10);
nor gn9_1_10(C1_10, n1_1_10, n5_1_10);

/* FA MFA2_10(S2_10,C2_10,S3_9,C2_9,A2B11); */
nor gn1_2_10(n1_2_10, S3_9, C2_9);
nor gn2_2_10(n2_2_10, n1_2_10, C2_9);
nor gn3_2_10(n3_2_10, S3_9, n1_2_10);
nor gn4_2_10(n4_2_10, n2_2_10, n3_2_10);
nor gn5_2_10(n5_2_10, A2B11, n4_2_10);
nor gn6_2_10(n6_2_10, A2B11, n5_2_10);
nor gn7_2_10(n7_2_10, n4_2_10, n5_2_10);
nor gn8_2_10(S2_10, n6_2_10, n7_2_10);
nor gn9_2_10(C2_10, n1_2_10, n5_2_10);

/* FA MFA3_10(S3_10,C3_10,S4_9,C3_9,A3B11); */
nor gn1_3_10(n1_3_10, S4_9, C3_9);
nor gn2_3_10(n2_3_10, n1_3_10, C3_9);
nor gn3_3_10(n3_3_10, S4_9, n1_3_10);
nor gn4_3_10(n4_3_10, n2_3_10, n3_3_10);
nor gn5_3_10(n5_3_10, A3B11, n4_3_10);
nor gn6_3_10(n6_3_10, A3B11, n5_3_10);
nor gn7_3_10(n7_3_10, n4_3_10, n5_3_10);
nor gn8_3_10(S3_10, n6_3_10, n7_3_10);
nor gn9_3_10(C3_10, n1_3_10, n5_3_10);

/* FA MFA4_10(S4_10,C4_10,S5_9,C4_9,A4B11); */
nor gn1_4_10(n1_4_10, S5_9, C4_9);
nor gn2_4_10(n2_4_10, n1_4_10, C4_9);
nor gn3_4_10(n3_4_10, S5_9, n1_4_10);
nor gn4_4_10(n4_4_10, n2_4_10, n3_4_10);
nor gn5_4_10(n5_4_10, A4B11, n4_4_10);
nor gn6_4_10(n6_4_10, A4B11, n5_4_10);
nor gn7_4_10(n7_4_10, n4_4_10, n5_4_10);
nor gn8_4_10(S4_10, n6_4_10, n7_4_10);
nor gn9_4_10(C4_10, n1_4_10, n5_4_10);

/* FA MFA5_10(S5_10,C5_10,S6_9,C5_9,A5B11); */
nor gn1_5_10(n1_5_10, S6_9, C5_9);
nor gn2_5_10(n2_5_10, n1_5_10, C5_9);
nor gn3_5_10(n3_5_10, S6_9, n1_5_10);
nor gn4_5_10(n4_5_10, n2_5_10, n3_5_10);
nor gn5_5_10(n5_5_10, A5B11, n4_5_10);
nor gn6_5_10(n6_5_10, A5B11, n5_5_10);
nor gn7_5_10(n7_5_10, n4_5_10, n5_5_10);
nor gn8_5_10(S5_10, n6_5_10, n7_5_10);
nor gn9_5_10(C5_10, n1_5_10, n5_5_10);

/* FA MFA6_10(S6_10,C6_10,S7_9,C6_9,A6B11); */
nor gn1_6_10(n1_6_10, S7_9, C6_9);
nor gn2_6_10(n2_6_10, n1_6_10, C6_9);
nor gn3_6_10(n3_6_10, S7_9, n1_6_10);
nor gn4_6_10(n4_6_10, n2_6_10, n3_6_10);
nor gn5_6_10(n5_6_10, A6B11, n4_6_10);
nor gn6_6_10(n6_6_10, A6B11, n5_6_10);
nor gn7_6_10(n7_6_10, n4_6_10, n5_6_10);
nor gn8_6_10(S6_10, n6_6_10, n7_6_10);
nor gn9_6_10(C6_10, n1_6_10, n5_6_10);

/* FA MFA7_10(S7_10,C7_10,S8_9,C7_9,A7B11); */
nor gn1_7_10(n1_7_10, S8_9, C7_9);
nor gn2_7_10(n2_7_10, n1_7_10, C7_9);
nor gn3_7_10(n3_7_10, S8_9, n1_7_10);
nor gn4_7_10(n4_7_10, n2_7_10, n3_7_10);
nor gn5_7_10(n5_7_10, A7B11, n4_7_10);
nor gn6_7_10(n6_7_10, A7B11, n5_7_10);
nor gn7_7_10(n7_7_10, n4_7_10, n5_7_10);
nor gn8_7_10(S7_10, n6_7_10, n7_7_10);
nor gn9_7_10(C7_10, n1_7_10, n5_7_10);

/* FA MFA8_10(S8_10,C8_10,S9_9,C8_9,A8B11); */
nor gn1_8_10(n1_8_10, S9_9, C8_9);
nor gn2_8_10(n2_8_10, n1_8_10, C8_9);
nor gn3_8_10(n3_8_10, S9_9, n1_8_10);
nor gn4_8_10(n4_8_10, n2_8_10, n3_8_10);
nor gn5_8_10(n5_8_10, A8B11, n4_8_10);
nor gn6_8_10(n6_8_10, A8B11, n5_8_10);
nor gn7_8_10(n7_8_10, n4_8_10, n5_8_10);
nor gn8_8_10(S8_10, n6_8_10, n7_8_10);
nor gn9_8_10(C8_10, n1_8_10, n5_8_10);

/* FA MFA9_10(S9_10,C9_10,S10_9,C9_9,A9B11); */
nor gn1_9_10(n1_9_10, S10_9, C9_9);
nor gn2_9_10(n2_9_10, n1_9_10, C9_9);
nor gn3_9_10(n3_9_10, S10_9, n1_9_10);
nor gn4_9_10(n4_9_10, n2_9_10, n3_9_10);
nor gn5_9_10(n5_9_10, A9B11, n4_9_10);
nor gn6_9_10(n6_9_10, A9B11, n5_9_10);
nor gn7_9_10(n7_9_10, n4_9_10, n5_9_10);
nor gn8_9_10(S9_10, n6_9_10, n7_9_10);
nor gn9_9_10(C9_10, n1_9_10, n5_9_10);

/* FA MFA10_10(S10_10,C10_10,S11_9,C10_9,A10B11); */
nor gn1_10_10(n1_10_10, S11_9, C10_9);
nor gn2_10_10(n2_10_10, n1_10_10, C10_9);
nor gn3_10_10(n3_10_10, S11_9, n1_10_10);
nor gn4_10_10(n4_10_10, n2_10_10, n3_10_10);
nor gn5_10_10(n5_10_10, A10B11, n4_10_10);
nor gn6_10_10(n6_10_10, A10B11, n5_10_10);
nor gn7_10_10(n7_10_10, n4_10_10, n5_10_10);
nor gn8_10_10(S10_10, n6_10_10, n7_10_10);
nor gn9_10_10(C10_10, n1_10_10, n5_10_10);

/* FA MFA11_10(S11_10,C11_10,S12_9,C11_9,A11B11); */
nor gn1_11_10(n1_11_10, S12_9, C11_9);
nor gn2_11_10(n2_11_10, n1_11_10, C11_9);
nor gn3_11_10(n3_11_10, S12_9, n1_11_10);
nor gn4_11_10(n4_11_10, n2_11_10, n3_11_10);
nor gn5_11_10(n5_11_10, A11B11, n4_11_10);
nor gn6_11_10(n6_11_10, A11B11, n5_11_10);
nor gn7_11_10(n7_11_10, n4_11_10, n5_11_10);
nor gn8_11_10(S11_10, n6_11_10, n7_11_10);
nor gn9_11_10(C11_10, n1_11_10, n5_11_10);

/* FA MFA12_10(S12_10,C12_10,S13_9,C12_9,A12B11); */
nor gn1_12_10(n1_12_10, S13_9, C12_9);
nor gn2_12_10(n2_12_10, n1_12_10, C12_9);
nor gn3_12_10(n3_12_10, S13_9, n1_12_10);
nor gn4_12_10(n4_12_10, n2_12_10, n3_12_10);
nor gn5_12_10(n5_12_10, A12B11, n4_12_10);
nor gn6_12_10(n6_12_10, A12B11, n5_12_10);
nor gn7_12_10(n7_12_10, n4_12_10, n5_12_10);
nor gn8_12_10(S12_10, n6_12_10, n7_12_10);
nor gn9_12_10(C12_10, n1_12_10, n5_12_10);

/* FA MFA13_10(S13_10,C13_10,S14_9,C13_9,A13B11); */
nor gn1_13_10(n1_13_10, S14_9, C13_9);
nor gn2_13_10(n2_13_10, n1_13_10, C13_9);
nor gn3_13_10(n3_13_10, S14_9, n1_13_10);
nor gn4_13_10(n4_13_10, n2_13_10, n3_13_10);
nor gn5_13_10(n5_13_10, A13B11, n4_13_10);
nor gn6_13_10(n6_13_10, A13B11, n5_13_10);
nor gn7_13_10(n7_13_10, n4_13_10, n5_13_10);
nor gn8_13_10(S13_10, n6_13_10, n7_13_10);
nor gn9_13_10(C13_10, n1_13_10, n5_13_10);

/* FA MFA14_10(S14_10,C14_10,A15B10,C14_9,A14B11); */
nor gn1_14_10(n1_14_10, A15B10, C14_9);
nor gn2_14_10(n2_14_10, n1_14_10, C14_9);
nor gn3_14_10(n3_14_10, A15B10, n1_14_10);
nor gn4_14_10(n4_14_10, n2_14_10, n3_14_10);
nor gn5_14_10(n5_14_10, A14B11, n4_14_10);
nor gn6_14_10(n6_14_10, A14B11, n5_14_10);
nor gn7_14_10(n7_14_10, n4_14_10, n5_14_10);
nor gn8_14_10(S14_10, n6_14_10, n7_14_10);
nor gn9_14_10(C14_10, n1_14_10, n5_14_10);

/* FA MFA0_11(S0_11,C0_11,S1_10,C0_10,A0B12); */
nor gn1_0_11(n1_0_11, S1_10, C0_10);
nor gn2_0_11(n2_0_11, n1_0_11, C0_10);
nor gn3_0_11(n3_0_11, S1_10, n1_0_11);
nor gn4_0_11(n4_0_11, n2_0_11, n3_0_11);
nor gn5_0_11(n5_0_11, A0B12, n4_0_11);
nor gn6_0_11(n6_0_11, A0B12, n5_0_11);
nor gn7_0_11(n7_0_11, n4_0_11, n5_0_11);
nor gn8_0_11(S0_11, n6_0_11, n7_0_11);
nor gn9_0_11(C0_11, n1_0_11, n5_0_11);

/* FA MFA1_11(S1_11,C1_11,S2_10,C1_10,A1B12); */
nor gn1_1_11(n1_1_11, S2_10, C1_10);
nor gn2_1_11(n2_1_11, n1_1_11, C1_10);
nor gn3_1_11(n3_1_11, S2_10, n1_1_11);
nor gn4_1_11(n4_1_11, n2_1_11, n3_1_11);
nor gn5_1_11(n5_1_11, A1B12, n4_1_11);
nor gn6_1_11(n6_1_11, A1B12, n5_1_11);
nor gn7_1_11(n7_1_11, n4_1_11, n5_1_11);
nor gn8_1_11(S1_11, n6_1_11, n7_1_11);
nor gn9_1_11(C1_11, n1_1_11, n5_1_11);

/* FA MFA2_11(S2_11,C2_11,S3_10,C2_10,A2B12); */
nor gn1_2_11(n1_2_11, S3_10, C2_10);
nor gn2_2_11(n2_2_11, n1_2_11, C2_10);
nor gn3_2_11(n3_2_11, S3_10, n1_2_11);
nor gn4_2_11(n4_2_11, n2_2_11, n3_2_11);
nor gn5_2_11(n5_2_11, A2B12, n4_2_11);
nor gn6_2_11(n6_2_11, A2B12, n5_2_11);
nor gn7_2_11(n7_2_11, n4_2_11, n5_2_11);
nor gn8_2_11(S2_11, n6_2_11, n7_2_11);
nor gn9_2_11(C2_11, n1_2_11, n5_2_11);

/* FA MFA3_11(S3_11,C3_11,S4_10,C3_10,A3B12); */
nor gn1_3_11(n1_3_11, S4_10, C3_10);
nor gn2_3_11(n2_3_11, n1_3_11, C3_10);
nor gn3_3_11(n3_3_11, S4_10, n1_3_11);
nor gn4_3_11(n4_3_11, n2_3_11, n3_3_11);
nor gn5_3_11(n5_3_11, A3B12, n4_3_11);
nor gn6_3_11(n6_3_11, A3B12, n5_3_11);
nor gn7_3_11(n7_3_11, n4_3_11, n5_3_11);
nor gn8_3_11(S3_11, n6_3_11, n7_3_11);
nor gn9_3_11(C3_11, n1_3_11, n5_3_11);

/* FA MFA4_11(S4_11,C4_11,S5_10,C4_10,A4B12); */
nor gn1_4_11(n1_4_11, S5_10, C4_10);
nor gn2_4_11(n2_4_11, n1_4_11, C4_10);
nor gn3_4_11(n3_4_11, S5_10, n1_4_11);
nor gn4_4_11(n4_4_11, n2_4_11, n3_4_11);
nor gn5_4_11(n5_4_11, A4B12, n4_4_11);
nor gn6_4_11(n6_4_11, A4B12, n5_4_11);
nor gn7_4_11(n7_4_11, n4_4_11, n5_4_11);
nor gn8_4_11(S4_11, n6_4_11, n7_4_11);
nor gn9_4_11(C4_11, n1_4_11, n5_4_11);

/* FA MFA5_11(S5_11,C5_11,S6_10,C5_10,A5B12); */
nor gn1_5_11(n1_5_11, S6_10, C5_10);
nor gn2_5_11(n2_5_11, n1_5_11, C5_10);
nor gn3_5_11(n3_5_11, S6_10, n1_5_11);
nor gn4_5_11(n4_5_11, n2_5_11, n3_5_11);
nor gn5_5_11(n5_5_11, A5B12, n4_5_11);
nor gn6_5_11(n6_5_11, A5B12, n5_5_11);
nor gn7_5_11(n7_5_11, n4_5_11, n5_5_11);
nor gn8_5_11(S5_11, n6_5_11, n7_5_11);
nor gn9_5_11(C5_11, n1_5_11, n5_5_11);

/* FA MFA6_11(S6_11,C6_11,S7_10,C6_10,A6B12); */
nor gn1_6_11(n1_6_11, S7_10, C6_10);
nor gn2_6_11(n2_6_11, n1_6_11, C6_10);
nor gn3_6_11(n3_6_11, S7_10, n1_6_11);
nor gn4_6_11(n4_6_11, n2_6_11, n3_6_11);
nor gn5_6_11(n5_6_11, A6B12, n4_6_11);
nor gn6_6_11(n6_6_11, A6B12, n5_6_11);
nor gn7_6_11(n7_6_11, n4_6_11, n5_6_11);
nor gn8_6_11(S6_11, n6_6_11, n7_6_11);
nor gn9_6_11(C6_11, n1_6_11, n5_6_11);

/* FA MFA7_11(S7_11,C7_11,S8_10,C7_10,A7B12); */
nor gn1_7_11(n1_7_11, S8_10, C7_10);
nor gn2_7_11(n2_7_11, n1_7_11, C7_10);
nor gn3_7_11(n3_7_11, S8_10, n1_7_11);
nor gn4_7_11(n4_7_11, n2_7_11, n3_7_11);
nor gn5_7_11(n5_7_11, A7B12, n4_7_11);
nor gn6_7_11(n6_7_11, A7B12, n5_7_11);
nor gn7_7_11(n7_7_11, n4_7_11, n5_7_11);
nor gn8_7_11(S7_11, n6_7_11, n7_7_11);
nor gn9_7_11(C7_11, n1_7_11, n5_7_11);

/* FA MFA8_11(S8_11,C8_11,S9_10,C8_10,A8B12); */
nor gn1_8_11(n1_8_11, S9_10, C8_10);
nor gn2_8_11(n2_8_11, n1_8_11, C8_10);
nor gn3_8_11(n3_8_11, S9_10, n1_8_11);
nor gn4_8_11(n4_8_11, n2_8_11, n3_8_11);
nor gn5_8_11(n5_8_11, A8B12, n4_8_11);
nor gn6_8_11(n6_8_11, A8B12, n5_8_11);
nor gn7_8_11(n7_8_11, n4_8_11, n5_8_11);
nor gn8_8_11(S8_11, n6_8_11, n7_8_11);
nor gn9_8_11(C8_11, n1_8_11, n5_8_11);

/* FA MFA9_11(S9_11,C9_11,S10_10,C9_10,A9B12); */
nor gn1_9_11(n1_9_11, S10_10, C9_10);
nor gn2_9_11(n2_9_11, n1_9_11, C9_10);
nor gn3_9_11(n3_9_11, S10_10, n1_9_11);
nor gn4_9_11(n4_9_11, n2_9_11, n3_9_11);
nor gn5_9_11(n5_9_11, A9B12, n4_9_11);
nor gn6_9_11(n6_9_11, A9B12, n5_9_11);
nor gn7_9_11(n7_9_11, n4_9_11, n5_9_11);
nor gn8_9_11(S9_11, n6_9_11, n7_9_11);
nor gn9_9_11(C9_11, n1_9_11, n5_9_11);

/* FA MFA10_11(S10_11,C10_11,S11_10,C10_10,A10B12); */
nor gn1_10_11(n1_10_11, S11_10, C10_10);
nor gn2_10_11(n2_10_11, n1_10_11, C10_10);
nor gn3_10_11(n3_10_11, S11_10, n1_10_11);
nor gn4_10_11(n4_10_11, n2_10_11, n3_10_11);
nor gn5_10_11(n5_10_11, A10B12, n4_10_11);
nor gn6_10_11(n6_10_11, A10B12, n5_10_11);
nor gn7_10_11(n7_10_11, n4_10_11, n5_10_11);
nor gn8_10_11(S10_11, n6_10_11, n7_10_11);
nor gn9_10_11(C10_11, n1_10_11, n5_10_11);

/* FA MFA11_11(S11_11,C11_11,S12_10,C11_10,A11B12); */
nor gn1_11_11(n1_11_11, S12_10, C11_10);
nor gn2_11_11(n2_11_11, n1_11_11, C11_10);
nor gn3_11_11(n3_11_11, S12_10, n1_11_11);
nor gn4_11_11(n4_11_11, n2_11_11, n3_11_11);
nor gn5_11_11(n5_11_11, A11B12, n4_11_11);
nor gn6_11_11(n6_11_11, A11B12, n5_11_11);
nor gn7_11_11(n7_11_11, n4_11_11, n5_11_11);
nor gn8_11_11(S11_11, n6_11_11, n7_11_11);
nor gn9_11_11(C11_11, n1_11_11, n5_11_11);

/* FA MFA12_11(S12_11,C12_11,S13_10,C12_10,A12B12); */
nor gn1_12_11(n1_12_11, S13_10, C12_10);
nor gn2_12_11(n2_12_11, n1_12_11, C12_10);
nor gn3_12_11(n3_12_11, S13_10, n1_12_11);
nor gn4_12_11(n4_12_11, n2_12_11, n3_12_11);
nor gn5_12_11(n5_12_11, A12B12, n4_12_11);
nor gn6_12_11(n6_12_11, A12B12, n5_12_11);
nor gn7_12_11(n7_12_11, n4_12_11, n5_12_11);
nor gn8_12_11(S12_11, n6_12_11, n7_12_11);
nor gn9_12_11(C12_11, n1_12_11, n5_12_11);

/* FA MFA13_11(S13_11,C13_11,S14_10,C13_10,A13B12); */
nor gn1_13_11(n1_13_11, S14_10, C13_10);
nor gn2_13_11(n2_13_11, n1_13_11, C13_10);
nor gn3_13_11(n3_13_11, S14_10, n1_13_11);
nor gn4_13_11(n4_13_11, n2_13_11, n3_13_11);
nor gn5_13_11(n5_13_11, A13B12, n4_13_11);
nor gn6_13_11(n6_13_11, A13B12, n5_13_11);
nor gn7_13_11(n7_13_11, n4_13_11, n5_13_11);
nor gn8_13_11(S13_11, n6_13_11, n7_13_11);
nor gn9_13_11(C13_11, n1_13_11, n5_13_11);

/* FA MFA14_11(S14_11,C14_11,A15B11,C14_10,A14B12); */
nor gn1_14_11(n1_14_11, A15B11, C14_10);
nor gn2_14_11(n2_14_11, n1_14_11, C14_10);
nor gn3_14_11(n3_14_11, A15B11, n1_14_11);
nor gn4_14_11(n4_14_11, n2_14_11, n3_14_11);
nor gn5_14_11(n5_14_11, A14B12, n4_14_11);
nor gn6_14_11(n6_14_11, A14B12, n5_14_11);
nor gn7_14_11(n7_14_11, n4_14_11, n5_14_11);
nor gn8_14_11(S14_11, n6_14_11, n7_14_11);
nor gn9_14_11(C14_11, n1_14_11, n5_14_11);

/* FA MFA0_12(S0_12,C0_12,S1_11,C0_11,A0B13); */
nor gn1_0_12(n1_0_12, S1_11, C0_11);
nor gn2_0_12(n2_0_12, n1_0_12, C0_11);
nor gn3_0_12(n3_0_12, S1_11, n1_0_12);
nor gn4_0_12(n4_0_12, n2_0_12, n3_0_12);
nor gn5_0_12(n5_0_12, A0B13, n4_0_12);
nor gn6_0_12(n6_0_12, A0B13, n5_0_12);
nor gn7_0_12(n7_0_12, n4_0_12, n5_0_12);
nor gn8_0_12(S0_12, n6_0_12, n7_0_12);
nor gn9_0_12(C0_12, n1_0_12, n5_0_12);

/* FA MFA1_12(S1_12,C1_12,S2_11,C1_11,A1B13); */
nor gn1_1_12(n1_1_12, S2_11, C1_11);
nor gn2_1_12(n2_1_12, n1_1_12, C1_11);
nor gn3_1_12(n3_1_12, S2_11, n1_1_12);
nor gn4_1_12(n4_1_12, n2_1_12, n3_1_12);
nor gn5_1_12(n5_1_12, A1B13, n4_1_12);
nor gn6_1_12(n6_1_12, A1B13, n5_1_12);
nor gn7_1_12(n7_1_12, n4_1_12, n5_1_12);
nor gn8_1_12(S1_12, n6_1_12, n7_1_12);
nor gn9_1_12(C1_12, n1_1_12, n5_1_12);

/* FA MFA2_12(S2_12,C2_12,S3_11,C2_11,A2B13); */
nor gn1_2_12(n1_2_12, S3_11, C2_11);
nor gn2_2_12(n2_2_12, n1_2_12, C2_11);
nor gn3_2_12(n3_2_12, S3_11, n1_2_12);
nor gn4_2_12(n4_2_12, n2_2_12, n3_2_12);
nor gn5_2_12(n5_2_12, A2B13, n4_2_12);
nor gn6_2_12(n6_2_12, A2B13, n5_2_12);
nor gn7_2_12(n7_2_12, n4_2_12, n5_2_12);
nor gn8_2_12(S2_12, n6_2_12, n7_2_12);
nor gn9_2_12(C2_12, n1_2_12, n5_2_12);

/* FA MFA3_12(S3_12,C3_12,S4_11,C3_11,A3B13); */
nor gn1_3_12(n1_3_12, S4_11, C3_11);
nor gn2_3_12(n2_3_12, n1_3_12, C3_11);
nor gn3_3_12(n3_3_12, S4_11, n1_3_12);
nor gn4_3_12(n4_3_12, n2_3_12, n3_3_12);
nor gn5_3_12(n5_3_12, A3B13, n4_3_12);
nor gn6_3_12(n6_3_12, A3B13, n5_3_12);
nor gn7_3_12(n7_3_12, n4_3_12, n5_3_12);
nor gn8_3_12(S3_12, n6_3_12, n7_3_12);
nor gn9_3_12(C3_12, n1_3_12, n5_3_12);

/* FA MFA4_12(S4_12,C4_12,S5_11,C4_11,A4B13); */
nor gn1_4_12(n1_4_12, S5_11, C4_11);
nor gn2_4_12(n2_4_12, n1_4_12, C4_11);
nor gn3_4_12(n3_4_12, S5_11, n1_4_12);
nor gn4_4_12(n4_4_12, n2_4_12, n3_4_12);
nor gn5_4_12(n5_4_12, A4B13, n4_4_12);
nor gn6_4_12(n6_4_12, A4B13, n5_4_12);
nor gn7_4_12(n7_4_12, n4_4_12, n5_4_12);
nor gn8_4_12(S4_12, n6_4_12, n7_4_12);
nor gn9_4_12(C4_12, n1_4_12, n5_4_12);

/* FA MFA5_12(S5_12,C5_12,S6_11,C5_11,A5B13); */
nor gn1_5_12(n1_5_12, S6_11, C5_11);
nor gn2_5_12(n2_5_12, n1_5_12, C5_11);
nor gn3_5_12(n3_5_12, S6_11, n1_5_12);
nor gn4_5_12(n4_5_12, n2_5_12, n3_5_12);
nor gn5_5_12(n5_5_12, A5B13, n4_5_12);
nor gn6_5_12(n6_5_12, A5B13, n5_5_12);
nor gn7_5_12(n7_5_12, n4_5_12, n5_5_12);
nor gn8_5_12(S5_12, n6_5_12, n7_5_12);
nor gn9_5_12(C5_12, n1_5_12, n5_5_12);

/* FA MFA6_12(S6_12,C6_12,S7_11,C6_11,A6B13); */
nor gn1_6_12(n1_6_12, S7_11, C6_11);
nor gn2_6_12(n2_6_12, n1_6_12, C6_11);
nor gn3_6_12(n3_6_12, S7_11, n1_6_12);
nor gn4_6_12(n4_6_12, n2_6_12, n3_6_12);
nor gn5_6_12(n5_6_12, A6B13, n4_6_12);
nor gn6_6_12(n6_6_12, A6B13, n5_6_12);
nor gn7_6_12(n7_6_12, n4_6_12, n5_6_12);
nor gn8_6_12(S6_12, n6_6_12, n7_6_12);
nor gn9_6_12(C6_12, n1_6_12, n5_6_12);

/* FA MFA7_12(S7_12,C7_12,S8_11,C7_11,A7B13); */
nor gn1_7_12(n1_7_12, S8_11, C7_11);
nor gn2_7_12(n2_7_12, n1_7_12, C7_11);
nor gn3_7_12(n3_7_12, S8_11, n1_7_12);
nor gn4_7_12(n4_7_12, n2_7_12, n3_7_12);
nor gn5_7_12(n5_7_12, A7B13, n4_7_12);
nor gn6_7_12(n6_7_12, A7B13, n5_7_12);
nor gn7_7_12(n7_7_12, n4_7_12, n5_7_12);
nor gn8_7_12(S7_12, n6_7_12, n7_7_12);
nor gn9_7_12(C7_12, n1_7_12, n5_7_12);

/* FA MFA8_12(S8_12,C8_12,S9_11,C8_11,A8B13); */
nor gn1_8_12(n1_8_12, S9_11, C8_11);
nor gn2_8_12(n2_8_12, n1_8_12, C8_11);
nor gn3_8_12(n3_8_12, S9_11, n1_8_12);
nor gn4_8_12(n4_8_12, n2_8_12, n3_8_12);
nor gn5_8_12(n5_8_12, A8B13, n4_8_12);
nor gn6_8_12(n6_8_12, A8B13, n5_8_12);
nor gn7_8_12(n7_8_12, n4_8_12, n5_8_12);
nor gn8_8_12(S8_12, n6_8_12, n7_8_12);
nor gn9_8_12(C8_12, n1_8_12, n5_8_12);

/* FA MFA9_12(S9_12,C9_12,S10_11,C9_11,A9B13); */
nor gn1_9_12(n1_9_12, S10_11, C9_11);
nor gn2_9_12(n2_9_12, n1_9_12, C9_11);
nor gn3_9_12(n3_9_12, S10_11, n1_9_12);
nor gn4_9_12(n4_9_12, n2_9_12, n3_9_12);
nor gn5_9_12(n5_9_12, A9B13, n4_9_12);
nor gn6_9_12(n6_9_12, A9B13, n5_9_12);
nor gn7_9_12(n7_9_12, n4_9_12, n5_9_12);
nor gn8_9_12(S9_12, n6_9_12, n7_9_12);
nor gn9_9_12(C9_12, n1_9_12, n5_9_12);

/* FA MFA10_12(S10_12,C10_12,S11_11,C10_11,A10B13); */
nor gn1_10_12(n1_10_12, S11_11, C10_11);
nor gn2_10_12(n2_10_12, n1_10_12, C10_11);
nor gn3_10_12(n3_10_12, S11_11, n1_10_12);
nor gn4_10_12(n4_10_12, n2_10_12, n3_10_12);
nor gn5_10_12(n5_10_12, A10B13, n4_10_12);
nor gn6_10_12(n6_10_12, A10B13, n5_10_12);
nor gn7_10_12(n7_10_12, n4_10_12, n5_10_12);
nor gn8_10_12(S10_12, n6_10_12, n7_10_12);
nor gn9_10_12(C10_12, n1_10_12, n5_10_12);

/* FA MFA11_12(S11_12,C11_12,S12_11,C11_11,A11B13); */
nor gn1_11_12(n1_11_12, S12_11, C11_11);
nor gn2_11_12(n2_11_12, n1_11_12, C11_11);
nor gn3_11_12(n3_11_12, S12_11, n1_11_12);
nor gn4_11_12(n4_11_12, n2_11_12, n3_11_12);
nor gn5_11_12(n5_11_12, A11B13, n4_11_12);
nor gn6_11_12(n6_11_12, A11B13, n5_11_12);
nor gn7_11_12(n7_11_12, n4_11_12, n5_11_12);
nor gn8_11_12(S11_12, n6_11_12, n7_11_12);
nor gn9_11_12(C11_12, n1_11_12, n5_11_12);

/* FA MFA12_12(S12_12,C12_12,S13_11,C12_11,A12B13); */
nor gn1_12_12(n1_12_12, S13_11, C12_11);
nor gn2_12_12(n2_12_12, n1_12_12, C12_11);
nor gn3_12_12(n3_12_12, S13_11, n1_12_12);
nor gn4_12_12(n4_12_12, n2_12_12, n3_12_12);
nor gn5_12_12(n5_12_12, A12B13, n4_12_12);
nor gn6_12_12(n6_12_12, A12B13, n5_12_12);
nor gn7_12_12(n7_12_12, n4_12_12, n5_12_12);
nor gn8_12_12(S12_12, n6_12_12, n7_12_12);
nor gn9_12_12(C12_12, n1_12_12, n5_12_12);

/* FA MFA13_12(S13_12,C13_12,S14_11,C13_11,A13B13); */
nor gn1_13_12(n1_13_12, S14_11, C13_11);
nor gn2_13_12(n2_13_12, n1_13_12, C13_11);
nor gn3_13_12(n3_13_12, S14_11, n1_13_12);
nor gn4_13_12(n4_13_12, n2_13_12, n3_13_12);
nor gn5_13_12(n5_13_12, A13B13, n4_13_12);
nor gn6_13_12(n6_13_12, A13B13, n5_13_12);
nor gn7_13_12(n7_13_12, n4_13_12, n5_13_12);
nor gn8_13_12(S13_12, n6_13_12, n7_13_12);
nor gn9_13_12(C13_12, n1_13_12, n5_13_12);

/* FA MFA14_12(S14_12,C14_12,A15B12,C14_11,A14B13); */
nor gn1_14_12(n1_14_12, A15B12, C14_11);
nor gn2_14_12(n2_14_12, n1_14_12, C14_11);
nor gn3_14_12(n3_14_12, A15B12, n1_14_12);
nor gn4_14_12(n4_14_12, n2_14_12, n3_14_12);
nor gn5_14_12(n5_14_12, A14B13, n4_14_12);
nor gn6_14_12(n6_14_12, A14B13, n5_14_12);
nor gn7_14_12(n7_14_12, n4_14_12, n5_14_12);
nor gn8_14_12(S14_12, n6_14_12, n7_14_12);
nor gn9_14_12(C14_12, n1_14_12, n5_14_12);

/* FA MFA0_13(S0_13,C0_13,S1_12,C0_12,A0B14); */
nor gn1_0_13(n1_0_13, S1_12, C0_12);
nor gn2_0_13(n2_0_13, n1_0_13, C0_12);
nor gn3_0_13(n3_0_13, S1_12, n1_0_13);
nor gn4_0_13(n4_0_13, n2_0_13, n3_0_13);
nor gn5_0_13(n5_0_13, A0B14, n4_0_13);
nor gn6_0_13(n6_0_13, A0B14, n5_0_13);
nor gn7_0_13(n7_0_13, n4_0_13, n5_0_13);
nor gn8_0_13(S0_13, n6_0_13, n7_0_13);
nor gn9_0_13(C0_13, n1_0_13, n5_0_13);

/* FA MFA1_13(S1_13,C1_13,S2_12,C1_12,A1B14); */
nor gn1_1_13(n1_1_13, S2_12, C1_12);
nor gn2_1_13(n2_1_13, n1_1_13, C1_12);
nor gn3_1_13(n3_1_13, S2_12, n1_1_13);
nor gn4_1_13(n4_1_13, n2_1_13, n3_1_13);
nor gn5_1_13(n5_1_13, A1B14, n4_1_13);
nor gn6_1_13(n6_1_13, A1B14, n5_1_13);
nor gn7_1_13(n7_1_13, n4_1_13, n5_1_13);
nor gn8_1_13(S1_13, n6_1_13, n7_1_13);
nor gn9_1_13(C1_13, n1_1_13, n5_1_13);

/* FA MFA2_13(S2_13,C2_13,S3_12,C2_12,A2B14); */
nor gn1_2_13(n1_2_13, S3_12, C2_12);
nor gn2_2_13(n2_2_13, n1_2_13, C2_12);
nor gn3_2_13(n3_2_13, S3_12, n1_2_13);
nor gn4_2_13(n4_2_13, n2_2_13, n3_2_13);
nor gn5_2_13(n5_2_13, A2B14, n4_2_13);
nor gn6_2_13(n6_2_13, A2B14, n5_2_13);
nor gn7_2_13(n7_2_13, n4_2_13, n5_2_13);
nor gn8_2_13(S2_13, n6_2_13, n7_2_13);
nor gn9_2_13(C2_13, n1_2_13, n5_2_13);

/* FA MFA3_13(S3_13,C3_13,S4_12,C3_12,A3B14); */
nor gn1_3_13(n1_3_13, S4_12, C3_12);
nor gn2_3_13(n2_3_13, n1_3_13, C3_12);
nor gn3_3_13(n3_3_13, S4_12, n1_3_13);
nor gn4_3_13(n4_3_13, n2_3_13, n3_3_13);
nor gn5_3_13(n5_3_13, A3B14, n4_3_13);
nor gn6_3_13(n6_3_13, A3B14, n5_3_13);
nor gn7_3_13(n7_3_13, n4_3_13, n5_3_13);
nor gn8_3_13(S3_13, n6_3_13, n7_3_13);
nor gn9_3_13(C3_13, n1_3_13, n5_3_13);

/* FA MFA4_13(S4_13,C4_13,S5_12,C4_12,A4B14); */
nor gn1_4_13(n1_4_13, S5_12, C4_12);
nor gn2_4_13(n2_4_13, n1_4_13, C4_12);
nor gn3_4_13(n3_4_13, S5_12, n1_4_13);
nor gn4_4_13(n4_4_13, n2_4_13, n3_4_13);
nor gn5_4_13(n5_4_13, A4B14, n4_4_13);
nor gn6_4_13(n6_4_13, A4B14, n5_4_13);
nor gn7_4_13(n7_4_13, n4_4_13, n5_4_13);
nor gn8_4_13(S4_13, n6_4_13, n7_4_13);
nor gn9_4_13(C4_13, n1_4_13, n5_4_13);

/* FA MFA5_13(S5_13,C5_13,S6_12,C5_12,A5B14); */
nor gn1_5_13(n1_5_13, S6_12, C5_12);
nor gn2_5_13(n2_5_13, n1_5_13, C5_12);
nor gn3_5_13(n3_5_13, S6_12, n1_5_13);
nor gn4_5_13(n4_5_13, n2_5_13, n3_5_13);
nor gn5_5_13(n5_5_13, A5B14, n4_5_13);
nor gn6_5_13(n6_5_13, A5B14, n5_5_13);
nor gn7_5_13(n7_5_13, n4_5_13, n5_5_13);
nor gn8_5_13(S5_13, n6_5_13, n7_5_13);
nor gn9_5_13(C5_13, n1_5_13, n5_5_13);

/* FA MFA6_13(S6_13,C6_13,S7_12,C6_12,A6B14); */
nor gn1_6_13(n1_6_13, S7_12, C6_12);
nor gn2_6_13(n2_6_13, n1_6_13, C6_12);
nor gn3_6_13(n3_6_13, S7_12, n1_6_13);
nor gn4_6_13(n4_6_13, n2_6_13, n3_6_13);
nor gn5_6_13(n5_6_13, A6B14, n4_6_13);
nor gn6_6_13(n6_6_13, A6B14, n5_6_13);
nor gn7_6_13(n7_6_13, n4_6_13, n5_6_13);
nor gn8_6_13(S6_13, n6_6_13, n7_6_13);
nor gn9_6_13(C6_13, n1_6_13, n5_6_13);

/* FA MFA7_13(S7_13,C7_13,S8_12,C7_12,A7B14); */
nor gn1_7_13(n1_7_13, S8_12, C7_12);
nor gn2_7_13(n2_7_13, n1_7_13, C7_12);
nor gn3_7_13(n3_7_13, S8_12, n1_7_13);
nor gn4_7_13(n4_7_13, n2_7_13, n3_7_13);
nor gn5_7_13(n5_7_13, A7B14, n4_7_13);
nor gn6_7_13(n6_7_13, A7B14, n5_7_13);
nor gn7_7_13(n7_7_13, n4_7_13, n5_7_13);
nor gn8_7_13(S7_13, n6_7_13, n7_7_13);
nor gn9_7_13(C7_13, n1_7_13, n5_7_13);

/* FA MFA8_13(S8_13,C8_13,S9_12,C8_12,A8B14); */
nor gn1_8_13(n1_8_13, S9_12, C8_12);
nor gn2_8_13(n2_8_13, n1_8_13, C8_12);
nor gn3_8_13(n3_8_13, S9_12, n1_8_13);
nor gn4_8_13(n4_8_13, n2_8_13, n3_8_13);
nor gn5_8_13(n5_8_13, A8B14, n4_8_13);
nor gn6_8_13(n6_8_13, A8B14, n5_8_13);
nor gn7_8_13(n7_8_13, n4_8_13, n5_8_13);
nor gn8_8_13(S8_13, n6_8_13, n7_8_13);
nor gn9_8_13(C8_13, n1_8_13, n5_8_13);

/* FA MFA9_13(S9_13,C9_13,S10_12,C9_12,A9B14); */
nor gn1_9_13(n1_9_13, S10_12, C9_12);
nor gn2_9_13(n2_9_13, n1_9_13, C9_12);
nor gn3_9_13(n3_9_13, S10_12, n1_9_13);
nor gn4_9_13(n4_9_13, n2_9_13, n3_9_13);
nor gn5_9_13(n5_9_13, A9B14, n4_9_13);
nor gn6_9_13(n6_9_13, A9B14, n5_9_13);
nor gn7_9_13(n7_9_13, n4_9_13, n5_9_13);
nor gn8_9_13(S9_13, n6_9_13, n7_9_13);
nor gn9_9_13(C9_13, n1_9_13, n5_9_13);

/* FA MFA10_13(S10_13,C10_13,S11_12,C10_12,A10B14); */
nor gn1_10_13(n1_10_13, S11_12, C10_12);
nor gn2_10_13(n2_10_13, n1_10_13, C10_12);
nor gn3_10_13(n3_10_13, S11_12, n1_10_13);
nor gn4_10_13(n4_10_13, n2_10_13, n3_10_13);
nor gn5_10_13(n5_10_13, A10B14, n4_10_13);
nor gn6_10_13(n6_10_13, A10B14, n5_10_13);
nor gn7_10_13(n7_10_13, n4_10_13, n5_10_13);
nor gn8_10_13(S10_13, n6_10_13, n7_10_13);
nor gn9_10_13(C10_13, n1_10_13, n5_10_13);

/* FA MFA11_13(S11_13,C11_13,S12_12,C11_12,A11B14); */
nor gn1_11_13(n1_11_13, S12_12, C11_12);
nor gn2_11_13(n2_11_13, n1_11_13, C11_12);
nor gn3_11_13(n3_11_13, S12_12, n1_11_13);
nor gn4_11_13(n4_11_13, n2_11_13, n3_11_13);
nor gn5_11_13(n5_11_13, A11B14, n4_11_13);
nor gn6_11_13(n6_11_13, A11B14, n5_11_13);
nor gn7_11_13(n7_11_13, n4_11_13, n5_11_13);
nor gn8_11_13(S11_13, n6_11_13, n7_11_13);
nor gn9_11_13(C11_13, n1_11_13, n5_11_13);

/* FA MFA12_13(S12_13,C12_13,S13_12,C12_12,A12B14); */
nor gn1_12_13(n1_12_13, S13_12, C12_12);
nor gn2_12_13(n2_12_13, n1_12_13, C12_12);
nor gn3_12_13(n3_12_13, S13_12, n1_12_13);
nor gn4_12_13(n4_12_13, n2_12_13, n3_12_13);
nor gn5_12_13(n5_12_13, A12B14, n4_12_13);
nor gn6_12_13(n6_12_13, A12B14, n5_12_13);
nor gn7_12_13(n7_12_13, n4_12_13, n5_12_13);
nor gn8_12_13(S12_13, n6_12_13, n7_12_13);
nor gn9_12_13(C12_13, n1_12_13, n5_12_13);

/* FA MFA13_13(S13_13,C13_13,S14_12,C13_12,A13B14); */
nor gn1_13_13(n1_13_13, S14_12, C13_12);
nor gn2_13_13(n2_13_13, n1_13_13, C13_12);
nor gn3_13_13(n3_13_13, S14_12, n1_13_13);
nor gn4_13_13(n4_13_13, n2_13_13, n3_13_13);
nor gn5_13_13(n5_13_13, A13B14, n4_13_13);
nor gn6_13_13(n6_13_13, A13B14, n5_13_13);
nor gn7_13_13(n7_13_13, n4_13_13, n5_13_13);
nor gn8_13_13(S13_13, n6_13_13, n7_13_13);
nor gn9_13_13(C13_13, n1_13_13, n5_13_13);

/* FA MFA14_13(S14_13,C14_13,A15B13,C14_12,A14B14); */
nor gn1_14_13(n1_14_13, A15B13, C14_12);
nor gn2_14_13(n2_14_13, n1_14_13, C14_12);
nor gn3_14_13(n3_14_13, A15B13, n1_14_13);
nor gn4_14_13(n4_14_13, n2_14_13, n3_14_13);
nor gn5_14_13(n5_14_13, A14B14, n4_14_13);
nor gn6_14_13(n6_14_13, A14B14, n5_14_13);
nor gn7_14_13(n7_14_13, n4_14_13, n5_14_13);
nor gn8_14_13(S14_13, n6_14_13, n7_14_13);
nor gn9_14_13(C14_13, n1_14_13, n5_14_13);

/* FA MFA0_14(S0_14,C0_14,S1_13,C0_13,A0B15); */
nor gn1_0_14(n1_0_14, S1_13, C0_13);
nor gn2_0_14(n2_0_14, n1_0_14, C0_13);
nor gn3_0_14(n3_0_14, S1_13, n1_0_14);
nor gn4_0_14(n4_0_14, n2_0_14, n3_0_14);
nor gn5_0_14(n5_0_14, A0B15, n4_0_14);
nor gn6_0_14(n6_0_14, A0B15, n5_0_14);
nor gn7_0_14(n7_0_14, n4_0_14, n5_0_14);
nor gn8_0_14(S0_14, n6_0_14, n7_0_14);
nor gn9_0_14(C0_14, n1_0_14, n5_0_14);

/* FA MFA1_14(S1_14,C1_14,S2_13,C1_13,A1B15); */
nor gn1_1_14(n1_1_14, S2_13, C1_13);
nor gn2_1_14(n2_1_14, n1_1_14, C1_13);
nor gn3_1_14(n3_1_14, S2_13, n1_1_14);
nor gn4_1_14(n4_1_14, n2_1_14, n3_1_14);
nor gn5_1_14(n5_1_14, A1B15, n4_1_14);
nor gn6_1_14(n6_1_14, A1B15, n5_1_14);
nor gn7_1_14(n7_1_14, n4_1_14, n5_1_14);
nor gn8_1_14(S1_14, n6_1_14, n7_1_14);
nor gn9_1_14(C1_14, n1_1_14, n5_1_14);

/* FA MFA2_14(S2_14,C2_14,S3_13,C2_13,A2B15); */
nor gn1_2_14(n1_2_14, S3_13, C2_13);
nor gn2_2_14(n2_2_14, n1_2_14, C2_13);
nor gn3_2_14(n3_2_14, S3_13, n1_2_14);
nor gn4_2_14(n4_2_14, n2_2_14, n3_2_14);
nor gn5_2_14(n5_2_14, A2B15, n4_2_14);
nor gn6_2_14(n6_2_14, A2B15, n5_2_14);
nor gn7_2_14(n7_2_14, n4_2_14, n5_2_14);
nor gn8_2_14(S2_14, n6_2_14, n7_2_14);
nor gn9_2_14(C2_14, n1_2_14, n5_2_14);

/* FA MFA3_14(S3_14,C3_14,S4_13,C3_13,A3B15); */
nor gn1_3_14(n1_3_14, S4_13, C3_13);
nor gn2_3_14(n2_3_14, n1_3_14, C3_13);
nor gn3_3_14(n3_3_14, S4_13, n1_3_14);
nor gn4_3_14(n4_3_14, n2_3_14, n3_3_14);
nor gn5_3_14(n5_3_14, A3B15, n4_3_14);
nor gn6_3_14(n6_3_14, A3B15, n5_3_14);
nor gn7_3_14(n7_3_14, n4_3_14, n5_3_14);
nor gn8_3_14(S3_14, n6_3_14, n7_3_14);
nor gn9_3_14(C3_14, n1_3_14, n5_3_14);

/* FA MFA4_14(S4_14,C4_14,S5_13,C4_13,A4B15); */
nor gn1_4_14(n1_4_14, S5_13, C4_13);
nor gn2_4_14(n2_4_14, n1_4_14, C4_13);
nor gn3_4_14(n3_4_14, S5_13, n1_4_14);
nor gn4_4_14(n4_4_14, n2_4_14, n3_4_14);
nor gn5_4_14(n5_4_14, A4B15, n4_4_14);
nor gn6_4_14(n6_4_14, A4B15, n5_4_14);
nor gn7_4_14(n7_4_14, n4_4_14, n5_4_14);
nor gn8_4_14(S4_14, n6_4_14, n7_4_14);
nor gn9_4_14(C4_14, n1_4_14, n5_4_14);

/* FA MFA5_14(S5_14,C5_14,S6_13,C5_13,A5B15); */
nor gn1_5_14(n1_5_14, S6_13, C5_13);
nor gn2_5_14(n2_5_14, n1_5_14, C5_13);
nor gn3_5_14(n3_5_14, S6_13, n1_5_14);
nor gn4_5_14(n4_5_14, n2_5_14, n3_5_14);
nor gn5_5_14(n5_5_14, A5B15, n4_5_14);
nor gn6_5_14(n6_5_14, A5B15, n5_5_14);
nor gn7_5_14(n7_5_14, n4_5_14, n5_5_14);
nor gn8_5_14(S5_14, n6_5_14, n7_5_14);
nor gn9_5_14(C5_14, n1_5_14, n5_5_14);

/* FA MFA6_14(S6_14,C6_14,S7_13,C6_13,A6B15); */
nor gn1_6_14(n1_6_14, S7_13, C6_13);
nor gn2_6_14(n2_6_14, n1_6_14, C6_13);
nor gn3_6_14(n3_6_14, S7_13, n1_6_14);
nor gn4_6_14(n4_6_14, n2_6_14, n3_6_14);
nor gn5_6_14(n5_6_14, A6B15, n4_6_14);
nor gn6_6_14(n6_6_14, A6B15, n5_6_14);
nor gn7_6_14(n7_6_14, n4_6_14, n5_6_14);
nor gn8_6_14(S6_14, n6_6_14, n7_6_14);
nor gn9_6_14(C6_14, n1_6_14, n5_6_14);

/* FA MFA7_14(S7_14,C7_14,S8_13,C7_13,A7B15); */
nor gn1_7_14(n1_7_14, S8_13, C7_13);
nor gn2_7_14(n2_7_14, n1_7_14, C7_13);
nor gn3_7_14(n3_7_14, S8_13, n1_7_14);
nor gn4_7_14(n4_7_14, n2_7_14, n3_7_14);
nor gn5_7_14(n5_7_14, A7B15, n4_7_14);
nor gn6_7_14(n6_7_14, A7B15, n5_7_14);
nor gn7_7_14(n7_7_14, n4_7_14, n5_7_14);
nor gn8_7_14(S7_14, n6_7_14, n7_7_14);
nor gn9_7_14(C7_14, n1_7_14, n5_7_14);

/* FA MFA8_14(S8_14,C8_14,S9_13,C8_13,A8B15); */
nor gn1_8_14(n1_8_14, S9_13, C8_13);
nor gn2_8_14(n2_8_14, n1_8_14, C8_13);
nor gn3_8_14(n3_8_14, S9_13, n1_8_14);
nor gn4_8_14(n4_8_14, n2_8_14, n3_8_14);
nor gn5_8_14(n5_8_14, A8B15, n4_8_14);
nor gn6_8_14(n6_8_14, A8B15, n5_8_14);
nor gn7_8_14(n7_8_14, n4_8_14, n5_8_14);
nor gn8_8_14(S8_14, n6_8_14, n7_8_14);
nor gn9_8_14(C8_14, n1_8_14, n5_8_14);

/* FA MFA9_14(S9_14,C9_14,S10_13,C9_13,A9B15); */
nor gn1_9_14(n1_9_14, S10_13, C9_13);
nor gn2_9_14(n2_9_14, n1_9_14, C9_13);
nor gn3_9_14(n3_9_14, S10_13, n1_9_14);
nor gn4_9_14(n4_9_14, n2_9_14, n3_9_14);
nor gn5_9_14(n5_9_14, A9B15, n4_9_14);
nor gn6_9_14(n6_9_14, A9B15, n5_9_14);
nor gn7_9_14(n7_9_14, n4_9_14, n5_9_14);
nor gn8_9_14(S9_14, n6_9_14, n7_9_14);
nor gn9_9_14(C9_14, n1_9_14, n5_9_14);

/* FA MFA10_14(S10_14,C10_14,S11_13,C10_13,A10B15); */
nor gn1_10_14(n1_10_14, S11_13, C10_13);
nor gn2_10_14(n2_10_14, n1_10_14, C10_13);
nor gn3_10_14(n3_10_14, S11_13, n1_10_14);
nor gn4_10_14(n4_10_14, n2_10_14, n3_10_14);
nor gn5_10_14(n5_10_14, A10B15, n4_10_14);
nor gn6_10_14(n6_10_14, A10B15, n5_10_14);
nor gn7_10_14(n7_10_14, n4_10_14, n5_10_14);
nor gn8_10_14(S10_14, n6_10_14, n7_10_14);
nor gn9_10_14(C10_14, n1_10_14, n5_10_14);

/* FA MFA11_14(S11_14,C11_14,S12_13,C11_13,A11B15); */
nor gn1_11_14(n1_11_14, S12_13, C11_13);
nor gn2_11_14(n2_11_14, n1_11_14, C11_13);
nor gn3_11_14(n3_11_14, S12_13, n1_11_14);
nor gn4_11_14(n4_11_14, n2_11_14, n3_11_14);
nor gn5_11_14(n5_11_14, A11B15, n4_11_14);
nor gn6_11_14(n6_11_14, A11B15, n5_11_14);
nor gn7_11_14(n7_11_14, n4_11_14, n5_11_14);
nor gn8_11_14(S11_14, n6_11_14, n7_11_14);
nor gn9_11_14(C11_14, n1_11_14, n5_11_14);

/* FA MFA12_14(S12_14,C12_14,S13_13,C12_13,A12B15); */
nor gn1_12_14(n1_12_14, S13_13, C12_13);
nor gn2_12_14(n2_12_14, n1_12_14, C12_13);
nor gn3_12_14(n3_12_14, S13_13, n1_12_14);
nor gn4_12_14(n4_12_14, n2_12_14, n3_12_14);
nor gn5_12_14(n5_12_14, A12B15, n4_12_14);
nor gn6_12_14(n6_12_14, A12B15, n5_12_14);
nor gn7_12_14(n7_12_14, n4_12_14, n5_12_14);
nor gn8_12_14(S12_14, n6_12_14, n7_12_14);
nor gn9_12_14(C12_14, n1_12_14, n5_12_14);

/* FA MFA13_14(S13_14,C13_14,S14_13,C13_13,A13B15); */
nor gn1_13_14(n1_13_14, S14_13, C13_13);
nor gn2_13_14(n2_13_14, n1_13_14, C13_13);
nor gn3_13_14(n3_13_14, S14_13, n1_13_14);
nor gn4_13_14(n4_13_14, n2_13_14, n3_13_14);
nor gn5_13_14(n5_13_14, A13B15, n4_13_14);
nor gn6_13_14(n6_13_14, A13B15, n5_13_14);
nor gn7_13_14(n7_13_14, n4_13_14, n5_13_14);
nor gn8_13_14(S13_14, n6_13_14, n7_13_14);
nor gn9_13_14(C13_14, n1_13_14, n5_13_14);

/* FA MFA14_14(S14_14,C14_14,A15B14,C14_13,A14B15); */
nor gn1_14_14(n1_14_14, A15B14, C14_13);
nor gn2_14_14(n2_14_14, n1_14_14, C14_13);
nor gn3_14_14(n3_14_14, A15B14, n1_14_14);
nor gn4_14_14(n4_14_14, n2_14_14, n3_14_14);
nor gn5_14_14(n5_14_14, A14B15, n4_14_14);
nor gn6_14_14(n6_14_14, A14B15, n5_14_14);
nor gn7_14_14(n7_14_14, n4_14_14, n5_14_14);
nor gn8_14_14(S14_14, n6_14_14, n7_14_14);
nor gn9_14_14(C14_14, n1_14_14, n5_14_14);

/* HA MHA0_15(S0_15,C0_15,S1_14,C0_14); */
nor gn1_0_15(n1_0_15, S1_14, C0_14);
nor gn2_0_15(n2_0_15, n1_0_15, C0_14);
nor gn3_0_15(n3_0_15, S1_14, n1_0_15);
nor gn4_0_15(n4_0_15, n2_0_15, n3_0_15);
not gn5_0_15(n5_0_15, n4_0_15);
not gn6_0_15(n6_0_15, n5_0_15);
nor gn7_0_15(n7_0_15, n4_0_15, n5_0_15);
nor gn8_0_15(S0_15, n6_0_15, n7_0_15);
nor gn9_0_15(C0_15, n1_0_15, n5_0_15);

/* FA MFA1_15(S1_15,C1_15,S2_14,C1_14,C0_15); */
nor gn1_1_15(n1_1_15, S2_14, C1_14);
nor gn2_1_15(n2_1_15, n1_1_15, C1_14);
nor gn3_1_15(n3_1_15, S2_14, n1_1_15);
nor gn4_1_15(n4_1_15, n2_1_15, n3_1_15);
nor gn5_1_15(n5_1_15, C0_15, n4_1_15);
nor gn6_1_15(n6_1_15, C0_15, n5_1_15);
nor gn7_1_15(n7_1_15, n4_1_15, n5_1_15);
nor gn8_1_15(S1_15, n6_1_15, n7_1_15);
nor gn9_1_15(C1_15, n1_1_15, n5_1_15);

/* FA MFA2_15(S2_15,C2_15,S3_14,C2_14,C1_15); */
nor gn1_2_15(n1_2_15, S3_14, C2_14);
nor gn2_2_15(n2_2_15, n1_2_15, C2_14);
nor gn3_2_15(n3_2_15, S3_14, n1_2_15);
nor gn4_2_15(n4_2_15, n2_2_15, n3_2_15);
nor gn5_2_15(n5_2_15, C1_15, n4_2_15);
nor gn6_2_15(n6_2_15, C1_15, n5_2_15);
nor gn7_2_15(n7_2_15, n4_2_15, n5_2_15);
nor gn8_2_15(S2_15, n6_2_15, n7_2_15);
nor gn9_2_15(C2_15, n1_2_15, n5_2_15);

/* FA MFA3_15(S3_15,C3_15,S4_14,C3_14,C2_15); */
nor gn1_3_15(n1_3_15, S4_14, C3_14);
nor gn2_3_15(n2_3_15, n1_3_15, C3_14);
nor gn3_3_15(n3_3_15, S4_14, n1_3_15);
nor gn4_3_15(n4_3_15, n2_3_15, n3_3_15);
nor gn5_3_15(n5_3_15, C2_15, n4_3_15);
nor gn6_3_15(n6_3_15, C2_15, n5_3_15);
nor gn7_3_15(n7_3_15, n4_3_15, n5_3_15);
nor gn8_3_15(S3_15, n6_3_15, n7_3_15);
nor gn9_3_15(C3_15, n1_3_15, n5_3_15);

/* FA MFA4_15(S4_15,C4_15,S5_14,C4_14,C3_15); */
nor gn1_4_15(n1_4_15, S5_14, C4_14);
nor gn2_4_15(n2_4_15, n1_4_15, C4_14);
nor gn3_4_15(n3_4_15, S5_14, n1_4_15);
nor gn4_4_15(n4_4_15, n2_4_15, n3_4_15);
nor gn5_4_15(n5_4_15, C3_15, n4_4_15);
nor gn6_4_15(n6_4_15, C3_15, n5_4_15);
nor gn7_4_15(n7_4_15, n4_4_15, n5_4_15);
nor gn8_4_15(S4_15, n6_4_15, n7_4_15);
nor gn9_4_15(C4_15, n1_4_15, n5_4_15);

/* FA MFA5_15(S5_15,C5_15,S6_14,C5_14,C4_15); */
nor gn1_5_15(n1_5_15, S6_14, C5_14);
nor gn2_5_15(n2_5_15, n1_5_15, C5_14);
nor gn3_5_15(n3_5_15, S6_14, n1_5_15);
nor gn4_5_15(n4_5_15, n2_5_15, n3_5_15);
nor gn5_5_15(n5_5_15, C4_15, n4_5_15);
nor gn6_5_15(n6_5_15, C4_15, n5_5_15);
nor gn7_5_15(n7_5_15, n4_5_15, n5_5_15);
nor gn8_5_15(S5_15, n6_5_15, n7_5_15);
nor gn9_5_15(C5_15, n1_5_15, n5_5_15);

/* FA MFA6_15(S6_15,C6_15,S7_14,C6_14,C5_15); */
nor gn1_6_15(n1_6_15, S7_14, C6_14);
nor gn2_6_15(n2_6_15, n1_6_15, C6_14);
nor gn3_6_15(n3_6_15, S7_14, n1_6_15);
nor gn4_6_15(n4_6_15, n2_6_15, n3_6_15);
nor gn5_6_15(n5_6_15, C5_15, n4_6_15);
nor gn6_6_15(n6_6_15, C5_15, n5_6_15);
nor gn7_6_15(n7_6_15, n4_6_15, n5_6_15);
nor gn8_6_15(S6_15, n6_6_15, n7_6_15);
nor gn9_6_15(C6_15, n1_6_15, n5_6_15);

/* FA MFA7_15(S7_15,C7_15,S8_14,C7_14,C6_15); */
nor gn1_7_15(n1_7_15, S8_14, C7_14);
nor gn2_7_15(n2_7_15, n1_7_15, C7_14);
nor gn3_7_15(n3_7_15, S8_14, n1_7_15);
nor gn4_7_15(n4_7_15, n2_7_15, n3_7_15);
nor gn5_7_15(n5_7_15, C6_15, n4_7_15);
nor gn6_7_15(n6_7_15, C6_15, n5_7_15);
nor gn7_7_15(n7_7_15, n4_7_15, n5_7_15);
nor gn8_7_15(S7_15, n6_7_15, n7_7_15);
nor gn9_7_15(C7_15, n1_7_15, n5_7_15);

/* FA MFA8_15(S8_15,C8_15,S9_14,C8_14,C7_15); */
nor gn1_8_15(n1_8_15, S9_14, C8_14);
nor gn2_8_15(n2_8_15, n1_8_15, C8_14);
nor gn3_8_15(n3_8_15, S9_14, n1_8_15);
nor gn4_8_15(n4_8_15, n2_8_15, n3_8_15);
nor gn5_8_15(n5_8_15, C7_15, n4_8_15);
nor gn6_8_15(n6_8_15, C7_15, n5_8_15);
nor gn7_8_15(n7_8_15, n4_8_15, n5_8_15);
nor gn8_8_15(S8_15, n6_8_15, n7_8_15);
nor gn9_8_15(C8_15, n1_8_15, n5_8_15);

/* FA MFA9_15(S9_15,C9_15,S10_14,C9_14,C8_15); */
nor gn1_9_15(n1_9_15, S10_14, C9_14);
nor gn2_9_15(n2_9_15, n1_9_15, C9_14);
nor gn3_9_15(n3_9_15, S10_14, n1_9_15);
nor gn4_9_15(n4_9_15, n2_9_15, n3_9_15);
nor gn5_9_15(n5_9_15, C8_15, n4_9_15);
nor gn6_9_15(n6_9_15, C8_15, n5_9_15);
nor gn7_9_15(n7_9_15, n4_9_15, n5_9_15);
nor gn8_9_15(S9_15, n6_9_15, n7_9_15);
nor gn9_9_15(C9_15, n1_9_15, n5_9_15);

/* FA MFA10_15(S10_15,C10_15,S11_14,C10_14,C9_15); */
nor gn1_10_15(n1_10_15, S11_14, C10_14);
nor gn2_10_15(n2_10_15, n1_10_15, C10_14);
nor gn3_10_15(n3_10_15, S11_14, n1_10_15);
nor gn4_10_15(n4_10_15, n2_10_15, n3_10_15);
nor gn5_10_15(n5_10_15, C9_15, n4_10_15);
nor gn6_10_15(n6_10_15, C9_15, n5_10_15);
nor gn7_10_15(n7_10_15, n4_10_15, n5_10_15);
nor gn8_10_15(S10_15, n6_10_15, n7_10_15);
nor gn9_10_15(C10_15, n1_10_15, n5_10_15);

/* FA MFA11_15(S11_15,C11_15,S12_14,C11_14,C10_15); */
nor gn1_11_15(n1_11_15, S12_14, C11_14);
nor gn2_11_15(n2_11_15, n1_11_15, C11_14);
nor gn3_11_15(n3_11_15, S12_14, n1_11_15);
nor gn4_11_15(n4_11_15, n2_11_15, n3_11_15);
nor gn5_11_15(n5_11_15, C10_15, n4_11_15);
nor gn6_11_15(n6_11_15, C10_15, n5_11_15);
nor gn7_11_15(n7_11_15, n4_11_15, n5_11_15);
nor gn8_11_15(S11_15, n6_11_15, n7_11_15);
nor gn9_11_15(C11_15, n1_11_15, n5_11_15);

/* FA MFA12_15(S12_15,C12_15,S13_14,C12_14,C11_15); */
nor gn1_12_15(n1_12_15, S13_14, C12_14);
nor gn2_12_15(n2_12_15, n1_12_15, C12_14);
nor gn3_12_15(n3_12_15, S13_14, n1_12_15);
nor gn4_12_15(n4_12_15, n2_12_15, n3_12_15);
nor gn5_12_15(n5_12_15, C11_15, n4_12_15);
nor gn6_12_15(n6_12_15, C11_15, n5_12_15);
nor gn7_12_15(n7_12_15, n4_12_15, n5_12_15);
nor gn8_12_15(S12_15, n6_12_15, n7_12_15);
nor gn9_12_15(C12_15, n1_12_15, n5_12_15);

/* FA MFA13_15(S13_15,C13_15,S14_14,C13_14,C12_15); */
nor gn1_13_15(n1_13_15, S14_14, C13_14);
nor gn2_13_15(n2_13_15, n1_13_15, C13_14);
nor gn3_13_15(n3_13_15, S14_14, n1_13_15);
nor gn4_13_15(n4_13_15, n2_13_15, n3_13_15);
nor gn5_13_15(n5_13_15, C12_15, n4_13_15);
nor gn6_13_15(n6_13_15, C12_15, n5_13_15);
nor gn7_13_15(n7_13_15, n4_13_15, n5_13_15);
nor gn8_13_15(S13_15, n6_13_15, n7_13_15);
nor gn9_13_15(C13_15, n1_13_15, n5_13_15);

/* FA MFA14_15(S14_15,C14_15,A15B15,C14_14,C13_15); */
nor gn1_14_15(n1_14_15, A15B15, C14_14);
nor gn2_14_15(n2_14_15, n1_14_15, C14_14);
nor gn3_14_15(n3_14_15, A15B15, n1_14_15);
nor gn4_14_15(n4_14_15, n2_14_15, n3_14_15);
nor gn5_14_15(n5_14_15, C13_15, n4_14_15);
nor gn6_14_15(n6_14_15, C13_15, n5_14_15);
nor gn7_14_15(n7_14_15, n4_14_15, n5_14_15);
nor gn8_14_15(S14_15, n6_14_15, n7_14_15);
nor gn9_14_15(C14_15, n1_14_15, n5_14_15);

endmodule /* TopLevel6288 */

/*************************************************************************/

